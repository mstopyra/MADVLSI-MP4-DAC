magic
tech sky130A
magscale 1 2
timestamp 1701223729
<< error_p >>
rect 7600 36400 9000 42400
rect 2000 29200 2200 35200
rect 7600 29200 7800 35200
rect 8800 29200 9000 35200
rect 14400 29200 14600 35200
rect 2800 21701 2801 27700
rect 4800 25400 5000 27700
rect 2800 21700 3000 21701
rect 6200 21700 6400 24200
rect 8200 21701 8201 27700
rect 11600 25400 11800 27700
rect 8200 21700 8400 21701
rect 10200 21700 10400 24200
rect 13600 21701 13601 27700
rect 13600 21700 13800 21701
rect 2800 14501 2801 20500
rect 6200 18000 6400 20500
rect 2800 14500 3000 14501
rect 4800 14500 5000 16800
rect 8200 14501 8201 20500
rect 10200 18000 10400 20500
rect 8200 14500 8400 14501
rect 11600 14500 11800 16800
rect 13600 14501 13601 20500
rect 13600 14500 13800 14501
rect 2000 7000 2200 13000
rect 7600 7000 7800 13000
rect 8800 7000 9000 13000
rect 14400 7000 14600 13000
rect 7600 -200 9000 5800
<< nwell >>
rect -2500 13500 19100 28300
<< nmos >>
rect -1000 36200 -200 42600
rect 2400 36200 3200 42600
rect 3800 36200 4600 42600
rect 6600 36200 7400 42600
rect 9200 36200 10000 42600
rect 12000 36200 12800 42600
rect 13400 36200 14200 42600
rect 16800 36200 17600 42600
rect -1000 29000 -200 35400
rect 2400 29000 3200 35400
rect 3800 29000 4600 35400
rect 6600 29000 7400 35400
rect 9200 29000 10000 35400
rect 12000 29000 12800 35400
rect 13400 29000 14200 35400
rect 16800 29000 17600 35400
rect -1000 6800 -200 13200
rect 2400 6800 3200 13200
rect 3800 6800 4600 13200
rect 6600 6800 7400 13200
rect 9200 6800 10000 13200
rect 12000 6800 12800 13200
rect 13400 6800 14200 13200
rect 16800 6800 17600 13200
rect -1000 -400 -200 6000
rect 2400 -400 3200 6000
rect 3800 -400 4600 6000
rect 6600 -400 7400 6000
rect 9200 -400 10000 6000
rect 12000 -400 12800 6000
rect 13400 -400 14200 6000
rect 16800 -400 17600 6000
<< pmos >>
rect 3800 21500 4600 27900
rect 5200 21500 6000 27900
rect 6600 21500 7400 27900
rect 9200 21500 10000 27900
rect 10600 21500 11400 27900
rect 12000 21500 12800 27900
rect 3800 14300 4600 20700
rect 5200 14300 6000 20700
rect 6600 14300 7400 20700
rect 9200 14300 10000 20700
rect 10600 14300 11400 20700
rect 12000 14300 12800 20700
<< ndiff >>
rect -1600 42400 -1000 42600
rect -1600 36400 -1400 42400
rect -1200 36400 -1000 42400
rect -1600 36200 -1000 36400
rect -200 42400 400 42600
rect -200 36400 0 42400
rect 200 36400 400 42400
rect -200 36200 400 36400
rect 1800 42400 2400 42600
rect 1800 36400 2000 42400
rect 2200 36400 2400 42400
rect 1800 36200 2400 36400
rect 3200 42400 3800 42600
rect 3200 36400 3400 42400
rect 3600 36400 3800 42400
rect 3200 36200 3800 36400
rect 4600 42400 5200 42600
rect 6000 42400 6600 42600
rect 4600 36400 4800 42400
rect 5000 36400 5200 42400
rect 6000 36400 6200 42400
rect 6400 36400 6600 42400
rect 4600 36200 5200 36400
rect 6000 36200 6600 36400
rect 7400 42400 9200 42600
rect 7400 36400 7600 42400
rect 9000 36400 9200 42400
rect 7400 36200 9200 36400
rect 10000 42400 10600 42600
rect 11400 42400 12000 42600
rect 10000 36400 10200 42400
rect 10400 36400 10600 42400
rect 11400 36400 11600 42400
rect 11800 36400 12000 42400
rect 10000 36200 10600 36400
rect 11400 36200 12000 36400
rect 12800 42400 13400 42600
rect 12800 36400 13000 42400
rect 13200 36400 13400 42400
rect 12800 36200 13400 36400
rect 14200 42400 14800 42600
rect 14200 36400 14400 42400
rect 14600 36400 14800 42400
rect 14200 36200 14800 36400
rect 16200 42400 16800 42600
rect 16200 36400 16400 42400
rect 16600 36400 16800 42400
rect 16200 36200 16800 36400
rect 17600 42400 18200 42600
rect 17600 36400 17800 42400
rect 18000 36400 18200 42400
rect 17600 36200 18200 36400
rect -1600 35200 -1000 35400
rect -1600 29200 -1400 35200
rect -1200 29200 -1000 35200
rect -1600 29000 -1000 29200
rect -200 35200 400 35400
rect -200 29200 0 35200
rect 200 29200 400 35200
rect -200 29000 400 29200
rect 1800 35200 2400 35400
rect 1800 29200 2000 35200
rect 2200 29200 2400 35200
rect 1800 29000 2400 29200
rect 3200 35200 3800 35400
rect 3200 29200 3400 35200
rect 3600 29200 3800 35200
rect 3200 29000 3800 29200
rect 4600 35200 5200 35400
rect 6000 35200 6600 35400
rect 4600 29200 4800 35200
rect 5000 29200 5200 35200
rect 6000 29200 6200 35200
rect 6400 29200 6600 35200
rect 4600 29000 5200 29200
rect 6000 29000 6600 29200
rect 7400 35200 8000 35400
rect 7400 29200 7600 35200
rect 7800 29200 8000 35200
rect 7400 29000 8000 29200
rect 8600 35200 9200 35400
rect 8600 29200 8800 35200
rect 9000 29200 9200 35200
rect 8600 29000 9200 29200
rect 10000 35200 10600 35400
rect 11400 35200 12000 35400
rect 10000 29200 10200 35200
rect 10400 29200 10600 35200
rect 11400 29200 11600 35200
rect 11800 29200 12000 35200
rect 10000 29000 10600 29200
rect 11400 29000 12000 29200
rect 12800 35200 13400 35400
rect 12800 29200 13000 35200
rect 13200 29200 13400 35200
rect 12800 29000 13400 29200
rect 14200 35200 14800 35400
rect 14200 29200 14400 35200
rect 14600 29200 14800 35200
rect 14200 29000 14800 29200
rect 16200 35200 16800 35400
rect 16200 29200 16400 35200
rect 16600 29200 16800 35200
rect 16200 29000 16800 29200
rect 17600 35200 18200 35400
rect 17600 29200 17800 35200
rect 18000 29200 18200 35200
rect 17600 29000 18200 29200
rect -1600 13000 -1000 13200
rect -1600 7000 -1400 13000
rect -1200 7000 -1000 13000
rect -1600 6800 -1000 7000
rect -200 13000 400 13200
rect -200 7000 0 13000
rect 200 7000 400 13000
rect -200 6800 400 7000
rect 1800 13000 2400 13200
rect 1800 7000 2000 13000
rect 2200 7000 2400 13000
rect 1800 6800 2400 7000
rect 3200 13000 3800 13200
rect 3200 7000 3400 13000
rect 3600 7000 3800 13000
rect 3200 6800 3800 7000
rect 4600 13000 5200 13200
rect 6000 13000 6600 13200
rect 4600 7000 4800 13000
rect 5000 7000 5200 13000
rect 6000 7000 6200 13000
rect 6400 7000 6600 13000
rect 4600 6800 5200 7000
rect 6000 6800 6600 7000
rect 7400 13000 8000 13200
rect 7400 7000 7600 13000
rect 7800 7000 8000 13000
rect 7400 6800 8000 7000
rect 8600 13000 9200 13200
rect 8600 7000 8800 13000
rect 9000 7000 9200 13000
rect 8600 6800 9200 7000
rect 10000 13000 10600 13200
rect 11400 13000 12000 13200
rect 10000 7000 10200 13000
rect 10400 7000 10600 13000
rect 11400 7000 11600 13000
rect 11800 7000 12000 13000
rect 10000 6800 10600 7000
rect 11400 6800 12000 7000
rect 12800 13000 13400 13200
rect 12800 7000 13000 13000
rect 13200 7000 13400 13000
rect 12800 6800 13400 7000
rect 14200 13000 14800 13200
rect 14200 7000 14400 13000
rect 14600 7000 14800 13000
rect 14200 6800 14800 7000
rect 16200 13000 16800 13200
rect 16200 7000 16400 13000
rect 16600 7000 16800 13000
rect 16200 6800 16800 7000
rect 17600 13000 18200 13200
rect 17600 7000 17800 13000
rect 18000 7000 18200 13000
rect 17600 6800 18200 7000
rect -1600 5800 -1000 6000
rect -1600 -200 -1400 5800
rect -1200 -200 -1000 5800
rect -1600 -400 -1000 -200
rect -200 5800 400 6000
rect -200 -200 0 5800
rect 200 -200 400 5800
rect -200 -400 400 -200
rect 1800 5800 2400 6000
rect 1800 -200 2000 5800
rect 2200 -200 2400 5800
rect 1800 -400 2400 -200
rect 3200 5800 3800 6000
rect 3200 -200 3400 5800
rect 3600 -200 3800 5800
rect 3200 -400 3800 -200
rect 4600 5800 5200 6000
rect 6000 5800 6600 6000
rect 4600 -200 4800 5800
rect 5000 -200 5200 5800
rect 6000 -200 6200 5800
rect 6400 -200 6600 5800
rect 4600 -400 5200 -200
rect 6000 -400 6600 -200
rect 7400 5800 9200 6000
rect 7400 -200 7600 5800
rect 9000 -200 9200 5800
rect 7400 -400 9200 -200
rect 10000 5800 10600 6000
rect 11400 5800 12000 6000
rect 10000 -200 10200 5800
rect 10400 -200 10600 5800
rect 11400 -200 11600 5800
rect 11800 -200 12000 5800
rect 10000 -400 10600 -200
rect 11400 -400 12000 -200
rect 12800 5800 13400 6000
rect 12800 -200 13000 5800
rect 13200 -200 13400 5800
rect 12800 -400 13400 -200
rect 14200 5800 14800 6000
rect 14200 -200 14400 5800
rect 14600 -200 14800 5800
rect 14200 -400 14800 -200
rect 16200 5800 16800 6000
rect 16200 -200 16400 5800
rect 16600 -200 16800 5800
rect 16200 -400 16800 -200
rect 17600 5800 18200 6000
rect 17600 -200 17800 5800
rect 18000 -200 18200 5800
rect 17600 -400 18200 -200
<< pdiff >>
rect 3200 27700 3800 27900
rect 3200 21700 3400 27700
rect 3600 21700 3800 27700
rect 3200 21500 3800 21700
rect 4600 27700 5200 27900
rect 4600 21700 4800 27700
rect 5000 21700 5200 27700
rect 4600 21500 5200 21700
rect 6000 27700 6600 27900
rect 6000 21700 6200 27700
rect 6400 21700 6600 27700
rect 6000 21500 6600 21700
rect 7400 27700 8000 27900
rect 8600 27700 9200 27900
rect 7400 21700 7600 27700
rect 7800 21700 8000 27700
rect 8600 21700 8800 27700
rect 9000 21700 9200 27700
rect 7400 21500 8000 21700
rect 8600 21500 9200 21700
rect 10000 27600 10600 27900
rect 10000 21700 10200 27600
rect 10400 21700 10600 27600
rect 10000 21500 10600 21700
rect 11400 27700 12000 27900
rect 11400 21700 11600 27700
rect 11800 21700 12000 27700
rect 11400 21500 12000 21700
rect 12800 27700 13400 27900
rect 12800 21700 13000 27700
rect 13200 21700 13400 27700
rect 12800 21500 13400 21700
rect 3200 20500 3800 20700
rect 3200 14500 3400 20500
rect 3600 14500 3800 20500
rect 3200 14300 3800 14500
rect 4600 20500 5200 20700
rect 4600 14500 4800 20500
rect 5000 14500 5200 20500
rect 4600 14300 5200 14500
rect 6000 20500 6600 20700
rect 6000 14500 6200 20500
rect 6400 14500 6600 20500
rect 6000 14300 6600 14500
rect 7400 20500 8000 20700
rect 8600 20500 9200 20700
rect 7400 14500 7600 20500
rect 7800 14500 8000 20500
rect 8600 14500 8800 20500
rect 9000 14500 9200 20500
rect 7400 14300 8000 14500
rect 8600 14300 9200 14500
rect 10000 20500 10600 20700
rect 10000 14500 10200 20500
rect 10400 14500 10600 20500
rect 10000 14300 10600 14500
rect 11400 20500 12000 20700
rect 11400 14500 11600 20500
rect 11800 14500 12000 20500
rect 11400 14300 12000 14500
rect 12800 20500 13400 20700
rect 12800 14500 13000 20500
rect 13200 14500 13400 20500
rect 12800 14300 13400 14500
<< ndiffc >>
rect -1400 36400 -1200 42400
rect 0 36400 200 42400
rect 2000 36400 2200 42400
rect 3400 36400 3600 42400
rect 4800 36400 5000 42400
rect 6200 36400 6400 42400
rect 7600 36400 9000 42400
rect 10200 36400 10400 42400
rect 11600 36400 11800 42400
rect 13000 36400 13200 42400
rect 14400 36400 14600 42400
rect 16400 36400 16600 42400
rect 17800 36400 18000 42400
rect -1400 29200 -1200 35200
rect 0 29200 200 35200
rect 2000 29200 2200 35200
rect 3400 29200 3600 35200
rect 4800 29200 5000 35200
rect 6200 29200 6400 35200
rect 7600 29200 7800 35200
rect 8800 29200 9000 35200
rect 10200 29200 10400 35200
rect 11600 29200 11800 35200
rect 13000 29200 13200 35200
rect 14400 29200 14600 35200
rect 16400 29200 16600 35200
rect 17800 29200 18000 35200
rect -1400 7000 -1200 13000
rect 0 7000 200 13000
rect 2000 7000 2200 13000
rect 3400 7000 3600 13000
rect 4800 7000 5000 13000
rect 6200 7000 6400 13000
rect 7600 7000 7800 13000
rect 8800 7000 9000 13000
rect 10200 7000 10400 13000
rect 11600 7000 11800 13000
rect 13000 7000 13200 13000
rect 14400 7000 14600 13000
rect 16400 7000 16600 13000
rect 17800 7000 18000 13000
rect -1400 -200 -1200 5800
rect 0 -200 200 5800
rect 2000 -200 2200 5800
rect 3400 -200 3600 5800
rect 4800 -200 5000 5800
rect 6200 -200 6400 5800
rect 7600 -200 9000 5800
rect 10200 -200 10400 5800
rect 11600 -200 11800 5800
rect 13000 -200 13200 5800
rect 14400 -200 14600 5800
rect 16400 -200 16600 5800
rect 17800 -200 18000 5800
<< pdiffc >>
rect 3400 21700 3600 27700
rect 4800 21700 5000 27700
rect 6200 21700 6400 27700
rect 7600 21700 7800 27700
rect 8800 21700 9000 27700
rect 10200 21700 10400 27600
rect 11600 21700 11800 27700
rect 13000 21700 13200 27700
rect 3400 14500 3600 20500
rect 4800 14500 5000 20500
rect 6200 14500 6400 20500
rect 7600 14500 7800 20500
rect 8800 14500 9000 20500
rect 10200 14500 10400 20500
rect 11600 14500 11800 20500
rect 13000 14500 13200 20500
<< psubdiff >>
rect -2400 42400 -1600 42600
rect -2400 36400 -2200 42400
rect -1800 36400 -1600 42400
rect -2400 36200 -1600 36400
rect 1000 42400 1800 42600
rect 1000 36400 1200 42400
rect 1600 36400 1800 42400
rect 1000 36200 1800 36400
rect 5200 42400 6000 42600
rect 5200 36400 5400 42400
rect 5800 36400 6000 42400
rect 5200 36200 6000 36400
rect 10600 42400 11400 42600
rect 10600 36400 10800 42400
rect 11200 36400 11400 42400
rect 10600 36200 11400 36400
rect 14800 42400 15600 42600
rect 14800 36400 15000 42400
rect 15400 36400 15600 42400
rect 14800 36200 15600 36400
rect 18200 42400 19000 42600
rect 18200 36400 18400 42400
rect 18800 36400 19000 42400
rect 18200 36200 19000 36400
rect -2400 35200 -1600 35400
rect -2400 29200 -2200 35200
rect -1800 29200 -1600 35200
rect -2400 29000 -1600 29200
rect 1000 35200 1800 35400
rect 1000 29200 1200 35200
rect 1600 29200 1800 35200
rect 1000 29000 1800 29200
rect 5200 35200 6000 35400
rect 5200 29200 5400 35200
rect 5800 29200 6000 35200
rect 5200 29000 6000 29200
rect 10600 35200 11400 35400
rect 10600 29200 10800 35200
rect 11200 29200 11400 35200
rect 10600 29000 11400 29200
rect 14800 35200 15600 35400
rect 14800 29200 15000 35200
rect 15400 29200 15600 35200
rect 14800 29000 15600 29200
rect 18200 35200 19000 35400
rect 18200 29200 18400 35200
rect 18800 29200 19000 35200
rect 18200 29000 19000 29200
rect -2400 13000 -1600 13200
rect -2400 7000 -2200 13000
rect -1800 7000 -1600 13000
rect -2400 6800 -1600 7000
rect 1000 13000 1800 13200
rect 1000 7000 1200 13000
rect 1600 7000 1800 13000
rect 1000 6800 1800 7000
rect 5200 13000 6000 13200
rect 5200 7000 5400 13000
rect 5800 7000 6000 13000
rect 5200 6800 6000 7000
rect 10600 13000 11400 13200
rect 10600 7000 10800 13000
rect 11200 7000 11400 13000
rect 10600 6800 11400 7000
rect 14800 13000 15600 13200
rect 14800 7000 15000 13000
rect 15400 7000 15600 13000
rect 14800 6800 15600 7000
rect 18200 13000 19000 13200
rect 18200 7000 18400 13000
rect 18800 7000 19000 13000
rect 18200 6800 19000 7000
rect -2400 5800 -1600 6000
rect -2400 -200 -2200 5800
rect -1800 -200 -1600 5800
rect -2400 -400 -1600 -200
rect 1000 5800 1800 6000
rect 1000 -200 1200 5800
rect 1600 -200 1800 5800
rect 1000 -400 1800 -200
rect 5200 5800 6000 6000
rect 5200 -200 5400 5800
rect 5800 -200 6000 5800
rect 5200 -400 6000 -200
rect 10600 5800 11400 6000
rect 10600 -200 10800 5800
rect 11200 -200 11400 5800
rect 10600 -400 11400 -200
rect 14800 5800 15600 6000
rect 14800 -200 15000 5800
rect 15400 -200 15600 5800
rect 14800 -400 15600 -200
rect 18200 5800 19000 6000
rect 18200 -200 18400 5800
rect 18800 -200 19000 5800
rect 18200 -400 19000 -200
<< nsubdiff >>
rect 2600 27700 3200 27900
rect 2600 21700 2800 27700
rect 3000 21700 3200 27700
rect 2600 21500 3200 21700
rect 8000 27700 8600 27900
rect 8000 21700 8200 27700
rect 8400 21700 8600 27700
rect 8000 21500 8600 21700
rect 13400 27700 14000 27900
rect 13400 21700 13600 27700
rect 13800 21700 14000 27700
rect 13400 21500 14000 21700
rect 2600 20500 3200 20700
rect 2600 14500 2800 20500
rect 3000 14500 3200 20500
rect 2600 14300 3200 14500
rect 8000 20500 8600 20700
rect 8000 14500 8200 20500
rect 8400 14500 8600 20500
rect 8000 14300 8600 14500
rect 13400 20500 14000 20700
rect 13400 14500 13600 20500
rect 13800 14500 14000 20500
rect 13400 14300 14000 14500
<< psubdiffcont >>
rect -2200 36400 -1800 42400
rect 1200 36400 1600 42400
rect 5400 36400 5800 42400
rect 10800 36400 11200 42400
rect 15000 36400 15400 42400
rect 18400 36400 18800 42400
rect -2200 29200 -1800 35200
rect 1200 29200 1600 35200
rect 5400 29200 5800 35200
rect 10800 29200 11200 35200
rect 15000 29200 15400 35200
rect 18400 29200 18800 35200
rect -2200 7000 -1800 13000
rect 1200 7000 1600 13000
rect 5400 7000 5800 13000
rect 10800 7000 11200 13000
rect 15000 7000 15400 13000
rect 18400 7000 18800 13000
rect -2200 -200 -1800 5800
rect 1200 -200 1600 5800
rect 5400 -200 5800 5800
rect 10800 -200 11200 5800
rect 15000 -200 15400 5800
rect 18400 -200 18800 5800
<< nsubdiffcont >>
rect 2800 21700 3000 27700
rect 8200 21700 8400 27700
rect 13600 21700 13800 27700
rect 2800 14500 3000 20500
rect 8200 14500 8400 20500
rect 13600 14500 13800 20500
<< poly >>
rect -1000 42600 -200 42800
rect 2400 42600 3200 42800
rect 3800 42600 4600 42800
rect 6600 42600 7400 42800
rect 9200 42600 10000 42800
rect 12000 42600 12800 42800
rect 13400 42600 14200 42800
rect 16800 42600 17600 42800
rect -1000 36100 -200 36200
rect -1000 35900 -900 36100
rect -300 35900 -200 36100
rect -1000 35800 -200 35900
rect -1000 35400 -200 35600
rect 2400 35400 3200 36200
rect 3800 35400 4600 36200
rect 6600 36000 7400 36200
rect 9200 36000 10000 36200
rect 6600 35900 10000 36000
rect 6600 35700 6700 35900
rect 9900 35700 10000 35900
rect 6600 35600 10000 35700
rect 6600 35400 7400 35500
rect 9200 35400 10000 35500
rect 12000 35400 12800 36200
rect 13400 35400 14200 36200
rect 16800 36100 17600 36200
rect 16800 35900 16900 36100
rect 17500 35900 17600 36100
rect 16800 35800 17600 35900
rect 16800 35400 17600 35600
rect -1000 28900 -200 29000
rect -1000 28700 -900 28900
rect -300 28700 -200 28900
rect -1000 28600 -200 28700
rect 2400 28900 3200 29000
rect 2400 28700 2500 28900
rect 3100 28700 3200 28900
rect 2400 28600 3200 28700
rect 3800 28900 4600 29000
rect 3800 28700 3900 28900
rect 4500 28700 4600 28900
rect 3800 28600 4600 28700
rect 6600 28800 7400 29000
rect 9200 28800 10000 29000
rect 6600 28700 10000 28800
rect 6600 28500 6700 28700
rect 9900 28500 10000 28700
rect 12000 28900 12800 29000
rect 12000 28700 12100 28900
rect 12700 28700 12800 28900
rect 12000 28600 12800 28700
rect 13400 28900 14200 29000
rect 13400 28700 13500 28900
rect 14100 28700 14200 28900
rect 13400 28600 14200 28700
rect 16800 28900 17600 29000
rect 16800 28700 16900 28900
rect 17500 28700 17600 28900
rect 16800 28600 17600 28700
rect 6600 28400 10000 28500
rect 3800 27900 4600 28000
rect 5200 27900 6000 28000
rect 6600 27900 7400 28000
rect 9200 27900 10000 28000
rect 10600 27900 11400 28000
rect 12000 27900 12800 28000
rect 3800 20700 4600 21500
rect 5200 21300 6000 21500
rect 6600 21300 7400 21500
rect 9200 21300 10000 21500
rect 10600 21300 11400 21500
rect 5200 21200 11400 21300
rect 5200 21000 6100 21200
rect 7300 21000 11400 21200
rect 5200 20900 11400 21000
rect 5200 20700 6000 20900
rect 6600 20700 7400 20900
rect 9200 20700 10000 20900
rect 10600 20700 11400 20900
rect 12000 20700 12800 21500
rect 3800 14200 4600 14300
rect 5200 14200 6000 14300
rect 6600 14200 7400 14300
rect 9200 14200 10000 14300
rect 10600 14200 11400 14300
rect 12000 14200 12800 14300
rect 3800 14000 3900 14200
rect 4500 14000 4600 14200
rect 3800 13900 4600 14000
rect 12000 14000 12100 14200
rect 12700 14000 12800 14200
rect 12000 13900 12800 14000
rect 6600 13700 10000 13800
rect -1000 13500 -200 13600
rect -1000 13300 -900 13500
rect -300 13300 -200 13500
rect -1000 13200 -200 13300
rect 2400 13500 3200 13600
rect 2400 13300 2500 13500
rect 3100 13300 3200 13500
rect 2400 13200 3200 13300
rect 3800 13500 4600 13600
rect 3800 13300 3900 13500
rect 4500 13300 4600 13500
rect 3800 13200 4600 13300
rect 6600 13500 6700 13700
rect 9900 13500 10000 13700
rect 6600 13400 10000 13500
rect 6600 13200 7400 13400
rect 9200 13200 10000 13400
rect 12000 13500 12800 13600
rect 12000 13300 12100 13500
rect 12700 13300 12800 13500
rect 12000 13200 12800 13300
rect 13400 13500 14200 13600
rect 13400 13300 13500 13500
rect 14100 13300 14200 13500
rect 13400 13200 14200 13300
rect 16800 13500 17600 13600
rect 16800 13300 16900 13500
rect 17500 13300 17600 13500
rect 16800 13200 17600 13300
rect -1000 6600 -200 6800
rect -1000 6300 -200 6400
rect -1000 6100 -900 6300
rect -300 6100 -200 6300
rect -1000 6000 -200 6100
rect 2400 6000 3200 6800
rect 3800 6000 4600 6800
rect 6600 6700 7400 6800
rect 9200 6700 10000 6800
rect 6600 6500 10000 6600
rect 6600 6300 6700 6500
rect 9900 6300 10000 6500
rect 6600 6200 10000 6300
rect 6600 6000 7400 6200
rect 9200 6000 10000 6200
rect 12000 6000 12800 6800
rect 13400 6000 14200 6800
rect 16800 6600 17600 6800
rect 16800 6300 17600 6400
rect 16800 6100 16900 6300
rect 17500 6100 17600 6300
rect 16800 6000 17600 6100
rect -1000 -600 -200 -400
rect 2400 -600 3200 -400
rect 3800 -600 4600 -400
rect 6600 -600 7400 -400
rect 9200 -600 10000 -400
rect 12000 -600 12800 -400
rect 13400 -600 14200 -400
rect 16800 -600 17600 -400
<< polycont >>
rect -900 35900 -300 36100
rect 6700 35700 9900 35900
rect 16900 35900 17500 36100
rect -900 28700 -300 28900
rect 2500 28700 3100 28900
rect 3900 28700 4500 28900
rect 6700 28500 9900 28700
rect 12100 28700 12700 28900
rect 13500 28700 14100 28900
rect 16900 28700 17500 28900
rect 6100 21000 7300 21200
rect 3900 14000 4500 14200
rect 12100 14000 12700 14200
rect -900 13300 -300 13500
rect 2500 13300 3100 13500
rect 3900 13300 4500 13500
rect 6700 13500 9900 13700
rect 12100 13300 12700 13500
rect 13500 13300 14100 13500
rect 16900 13300 17500 13500
rect -900 6100 -300 6300
rect 6700 6300 9900 6500
rect 16900 6100 17500 6300
<< locali >>
rect 1900 42600 5100 43000
rect -2300 42400 -1100 42500
rect -2300 36400 -2200 42400
rect -1800 36400 -1400 42400
rect -1200 36400 -1100 42400
rect -2300 36200 -1100 36400
rect -100 42400 300 42500
rect -100 36400 0 42400
rect 200 36400 300 42400
rect -2300 36100 -200 36200
rect -2300 35900 -900 36100
rect -300 35900 -200 36100
rect -2300 35800 -200 35900
rect -100 36000 300 36400
rect 1100 42400 1700 42500
rect 1100 36400 1200 42400
rect 1600 36400 1700 42400
rect 1100 36300 1700 36400
rect 1900 42400 2300 42600
rect 1900 36400 2000 42400
rect 2200 36400 2300 42400
rect 1900 36000 2300 36400
rect -2300 35200 -1100 35800
rect -2300 29200 -2200 35200
rect -1800 29200 -1400 35200
rect -1200 29200 -1100 35200
rect -2300 29000 -1100 29200
rect -100 35600 2300 36000
rect -100 35200 300 35600
rect -100 29200 0 35200
rect 200 29200 300 35200
rect -100 29000 300 29200
rect 1100 35200 1700 35300
rect 1100 29200 1200 35200
rect 1600 29200 1700 35200
rect 1100 29100 1700 29200
rect 1900 35200 2300 35600
rect 1900 29200 2000 35200
rect 2200 29200 2300 35200
rect 1900 29100 2300 29200
rect 3300 42400 3700 42500
rect 3300 36400 3400 42400
rect 3600 36400 3700 42400
rect 3300 35200 3700 36400
rect 3300 29200 3400 35200
rect 3600 29200 3700 35200
rect 3300 29000 3700 29200
rect 4700 42400 5100 42600
rect 11500 42600 14700 43000
rect 4700 36400 4800 42400
rect 5000 36400 5100 42400
rect 4700 36000 5100 36400
rect 5300 42400 5900 42500
rect 5300 36400 5400 42400
rect 5800 36400 5900 42400
rect 5300 36300 5900 36400
rect 6100 42400 6500 42500
rect 6100 36400 6200 42400
rect 6400 36400 6500 42400
rect 6100 36000 6500 36400
rect 7500 42400 9100 42500
rect 7500 36400 7600 42400
rect 9000 36400 9100 42400
rect 7500 36300 9100 36400
rect 10100 42400 10500 42500
rect 10100 36400 10200 42400
rect 10400 36400 10500 42400
rect 10100 36000 10500 36400
rect 10700 42400 11300 42500
rect 10700 36400 10800 42400
rect 11200 36400 11300 42400
rect 10700 36300 11300 36400
rect 11500 42400 11900 42600
rect 11500 36400 11600 42400
rect 11800 36400 11900 42400
rect 11500 36000 11900 36400
rect 12900 42400 13300 42500
rect 12900 36400 13000 42400
rect 13200 36400 13300 42400
rect 12900 36200 13300 36400
rect 14300 42400 14700 42600
rect 14300 36400 14400 42400
rect 14600 36400 14700 42400
rect 4700 35600 6500 36000
rect 6600 35900 10000 36000
rect 6600 35700 6700 35900
rect 9900 35700 10000 35900
rect 6600 35600 10000 35700
rect 10100 35600 11900 36000
rect 4700 35200 5100 35600
rect 4700 29200 4800 35200
rect 5000 29200 5100 35200
rect 4700 29100 5100 29200
rect 5300 35200 5900 35300
rect 5300 29200 5400 35200
rect 5800 29200 5900 35200
rect 5300 29100 5900 29200
rect 6100 35200 6500 35600
rect 6100 29200 6200 35200
rect 6400 29200 6500 35200
rect 6100 29100 6500 29200
rect 7500 35200 7900 35300
rect 7500 29200 7600 35200
rect 7800 29200 7900 35200
rect 7500 29100 7900 29200
rect 8700 35200 9100 35300
rect 8700 29200 8800 35200
rect 9000 29200 9100 35200
rect 10100 35200 10500 35600
rect 10100 29200 10200 35200
rect 10400 29200 10500 35200
rect 10700 35200 11300 35300
rect 10700 29200 10800 35200
rect 11200 29200 11300 35200
rect -2300 28900 -200 29000
rect -2300 28700 -900 28900
rect -300 28700 -200 28900
rect -2300 28600 -200 28700
rect 2400 28900 5100 29000
rect 2400 28700 2500 28900
rect 3100 28700 3900 28900
rect 4500 28700 5100 28900
rect 8700 28800 9100 29200
rect 10700 29100 11300 29200
rect 11500 35200 11900 35600
rect 12800 36100 13400 36200
rect 12800 35500 12900 36100
rect 13300 35500 13400 36100
rect 12800 35400 13400 35500
rect 14300 36000 14700 36400
rect 14900 42400 15500 42500
rect 14900 36400 15000 42400
rect 15400 36400 15500 42400
rect 14900 36300 15500 36400
rect 16300 42400 16700 42500
rect 16300 36400 16400 42400
rect 16600 36400 16700 42400
rect 16300 36000 16700 36400
rect 17700 42400 18900 42500
rect 17700 36400 17800 42400
rect 18000 36400 18400 42400
rect 18800 36400 18900 42400
rect 17700 36200 18900 36400
rect 14300 35600 16700 36000
rect 16800 36100 18900 36200
rect 16800 35900 16900 36100
rect 17500 35900 18900 36100
rect 16800 35800 18900 35900
rect 11500 29200 11600 35200
rect 11800 29200 11900 35200
rect 11500 29100 11900 29200
rect 12900 35200 13300 35400
rect 12900 29200 13000 35200
rect 13200 29200 13300 35200
rect 12900 29000 13300 29200
rect 14300 35200 14700 35600
rect 14300 29200 14400 35200
rect 14600 29200 14700 35200
rect 14300 29100 14700 29200
rect 14900 35200 15500 35300
rect 14900 29200 15000 35200
rect 15400 29200 15500 35200
rect 14900 29100 15500 29200
rect 16300 35200 16700 35600
rect 16300 29200 16400 35200
rect 16600 29200 16700 35200
rect 16300 29100 16700 29200
rect 17700 35200 18900 35800
rect 17700 29200 17800 35200
rect 18000 29200 18400 35200
rect 18800 29200 18900 35200
rect 17700 29000 18900 29200
rect 11500 28900 14200 29000
rect 2400 28600 5100 28700
rect 2700 27700 3700 27800
rect 2700 21700 2800 27700
rect 3000 21700 3400 27700
rect 3600 21700 3700 27700
rect 2700 21600 3700 21700
rect 4700 27700 5100 28600
rect 6600 28700 10000 28800
rect 6600 28500 6700 28700
rect 9900 28500 10000 28700
rect 6600 28400 10000 28500
rect 11500 28700 12100 28900
rect 12700 28700 13500 28900
rect 14100 28700 14200 28900
rect 11500 28600 14200 28700
rect 16800 28900 18900 29000
rect 16800 28700 16900 28900
rect 17500 28700 18900 28900
rect 16800 28600 18900 28700
rect 4700 21700 4800 27700
rect 5000 21700 5100 27700
rect 4700 21600 5100 21700
rect 6100 27700 6500 27800
rect 6100 21700 6200 27700
rect 6400 21700 6500 27700
rect 6100 21600 6500 21700
rect 7500 27700 9100 27800
rect 11500 27700 11900 28600
rect 7500 21700 7600 27700
rect 7800 21700 8200 27700
rect 8400 21700 8800 27700
rect 9000 21700 9100 27700
rect 7500 21600 9100 21700
rect 10100 27600 10500 27700
rect 10100 21700 10200 27600
rect 10400 21700 10500 27600
rect 10100 21600 10500 21700
rect 11500 21700 11600 27700
rect 11800 21700 11900 27700
rect 11500 21600 11900 21700
rect 12900 27700 13900 27800
rect 12900 21700 13000 27700
rect 13200 21700 13600 27700
rect 13800 21700 13900 27700
rect 12900 21600 13900 21700
rect 6000 21200 7400 21300
rect 6000 21000 6100 21200
rect 7300 21000 7400 21200
rect 6000 20900 7400 21000
rect 2700 20500 3700 20600
rect 2700 14500 2800 20500
rect 3000 14500 3400 20500
rect 3600 14500 3700 20500
rect 2700 14400 3700 14500
rect 4700 20500 5100 20600
rect 4700 14500 4800 20500
rect 5000 14500 5100 20500
rect 3800 14200 4600 14300
rect 3800 14000 3900 14200
rect 4500 14000 4600 14200
rect 3800 13900 4600 14000
rect 4700 13600 5100 14500
rect 6100 20500 6500 20600
rect 6100 14500 6200 20500
rect 6400 14500 6500 20500
rect 6100 14400 6500 14500
rect 7500 20500 9100 20600
rect 7500 14500 7600 20500
rect 7800 14500 8200 20500
rect 8400 14500 8800 20500
rect 9000 14500 9100 20500
rect 7500 14400 9100 14500
rect 10100 20500 10500 20600
rect 10100 14500 10200 20500
rect 10400 14500 10500 20500
rect 10100 14400 10500 14500
rect 11500 20500 11900 20600
rect 11500 14500 11600 20500
rect 11800 14500 11900 20500
rect -2300 13500 -200 13600
rect -2300 13300 -900 13500
rect -300 13300 -200 13500
rect -2300 13200 -200 13300
rect 2400 13500 5100 13600
rect 2400 13300 2500 13500
rect 3100 13300 3900 13500
rect 4500 13300 5100 13500
rect 6600 13700 10000 13800
rect 6600 13500 6700 13700
rect 9900 13500 10000 13700
rect 6600 13400 10000 13500
rect 11500 13600 11900 14500
rect 12900 20500 13900 20600
rect 12900 14500 13000 20500
rect 13200 14500 13600 20500
rect 13800 14500 13900 20500
rect 12900 14400 13900 14500
rect 12000 14200 12800 14300
rect 12000 14000 12100 14200
rect 12700 14000 12800 14200
rect 12000 13900 12800 14000
rect 18300 13600 18900 28600
rect 11500 13500 14200 13600
rect 2400 13200 5100 13300
rect -2300 13000 -1100 13200
rect -2300 7000 -2200 13000
rect -1800 7000 -1400 13000
rect -1200 7000 -1100 13000
rect -2300 6400 -1100 7000
rect -100 13000 300 13100
rect -100 7000 0 13000
rect 200 7000 300 13000
rect -100 6600 300 7000
rect 1100 13000 1700 13100
rect 1100 7000 1200 13000
rect 1600 7000 1700 13000
rect 1100 6900 1700 7000
rect 1900 13000 2300 13100
rect 1900 7000 2000 13000
rect 2200 7000 2300 13000
rect 1900 6600 2300 7000
rect 3300 13000 3700 13200
rect 3300 7000 3400 13000
rect 3600 7000 3700 13000
rect 3300 6800 3700 7000
rect 4700 13000 5100 13100
rect 4700 7000 4800 13000
rect 5000 7000 5100 13000
rect -2300 6300 -200 6400
rect -2300 6100 -900 6300
rect -300 6100 -200 6300
rect -2300 6000 -200 6100
rect -100 6200 2300 6600
rect -2300 5800 -1100 6000
rect -2300 -200 -2200 5800
rect -1800 -200 -1400 5800
rect -1200 -200 -1100 5800
rect -2300 -300 -1100 -200
rect -100 5800 300 6200
rect -100 -200 0 5800
rect 200 -200 300 5800
rect -100 -300 300 -200
rect 1100 5800 1700 5900
rect 1100 -200 1200 5800
rect 1600 -200 1700 5800
rect 1100 -300 1700 -200
rect 1900 5800 2300 6200
rect 3200 6700 3800 6800
rect 3200 6100 3300 6700
rect 3700 6100 3800 6700
rect 3200 6000 3800 6100
rect 4700 6600 5100 7000
rect 5300 13000 5900 13100
rect 7500 13000 7900 13400
rect 11500 13300 12100 13500
rect 12700 13300 13500 13500
rect 14100 13300 14200 13500
rect 11500 13200 14200 13300
rect 16800 13500 18900 13600
rect 16800 13300 16900 13500
rect 17500 13300 18900 13500
rect 16800 13200 18900 13300
rect 5300 7000 5400 13000
rect 5800 7000 5900 13000
rect 5300 6900 5900 7000
rect 6100 7000 6200 13000
rect 6400 7000 6500 13000
rect 6100 6600 6500 7000
rect 7500 7000 7600 13000
rect 7800 7000 7900 13000
rect 7500 6900 7900 7000
rect 8700 13000 9100 13100
rect 8700 7000 8800 13000
rect 9000 7000 9100 13000
rect 8700 6900 9100 7000
rect 10100 13000 10500 13100
rect 10100 7000 10200 13000
rect 10400 7000 10500 13000
rect 10100 6600 10500 7000
rect 10700 13000 11300 13100
rect 10700 7000 10800 13000
rect 11200 7000 11300 13000
rect 10700 6900 11300 7000
rect 11500 13000 11900 13100
rect 11500 7000 11600 13000
rect 11800 7000 11900 13000
rect 11500 6600 11900 7000
rect 4700 6200 6500 6600
rect 6600 6500 10000 6600
rect 6600 6300 6700 6500
rect 9900 6300 10000 6500
rect 6600 6200 10000 6300
rect 10100 6200 11900 6600
rect 1900 -200 2000 5800
rect 2200 -200 2300 5800
rect 1900 -400 2300 -200
rect 3300 5800 3700 6000
rect 3300 -200 3400 5800
rect 3600 -200 3700 5800
rect 3300 -300 3700 -200
rect 4700 5800 5100 6200
rect 4700 -200 4800 5800
rect 5000 -200 5100 5800
rect 4700 -400 5100 -200
rect 5300 5800 5900 5900
rect 5300 -200 5400 5800
rect 5800 -200 5900 5800
rect 5300 -300 5900 -200
rect 6100 5800 6500 6200
rect 6100 -200 6200 5800
rect 6400 -200 6500 5800
rect 6100 -300 6500 -200
rect 7500 5800 9100 5900
rect 7500 -200 7600 5800
rect 9000 -200 9100 5800
rect 7500 -300 9100 -200
rect 10100 5800 10500 6200
rect 10100 -200 10200 5800
rect 10400 -200 10500 5800
rect 10100 -300 10500 -200
rect 10700 5800 11300 5900
rect 10700 -200 10800 5800
rect 11200 -200 11300 5800
rect 10700 -300 11300 -200
rect 11500 5800 11900 6200
rect 11500 -200 11600 5800
rect 11800 -200 11900 5800
rect 11500 -300 11900 -200
rect 12900 13000 13300 13200
rect 12900 7000 13000 13000
rect 13200 7000 13300 13000
rect 12900 5800 13300 7000
rect 12900 -200 13000 5800
rect 13200 -200 13300 5800
rect 12900 -300 13300 -200
rect 14300 13000 14700 13100
rect 14300 7000 14400 13000
rect 14600 7000 14700 13000
rect 14300 6600 14700 7000
rect 14900 13000 15500 13100
rect 14900 7000 15000 13000
rect 15400 7000 15500 13000
rect 14900 6900 15500 7000
rect 16300 13000 16700 13200
rect 16300 7000 16400 13000
rect 16600 7000 16700 13000
rect 16300 6600 16700 7000
rect 14300 6200 16700 6600
rect 17700 13000 18900 13200
rect 17700 7000 17800 13000
rect 18000 7000 18400 13000
rect 18800 7000 18900 13000
rect 17700 6400 18900 7000
rect 14300 5800 14700 6200
rect 14300 -200 14400 5800
rect 14600 -200 14700 5800
rect 14300 -300 14700 -200
rect 14900 5800 15500 5900
rect 14900 -200 15000 5800
rect 15400 -200 15500 5800
rect 14900 -300 15500 -200
rect 16300 5800 16700 6200
rect 16800 6300 18900 6400
rect 16800 6100 16900 6300
rect 17500 6100 18900 6300
rect 16800 6000 18900 6100
rect 16300 -200 16400 5800
rect 16600 -200 16700 5800
rect 16300 -300 16700 -200
rect 17700 5800 18900 6000
rect 17700 -200 17800 5800
rect 18000 -200 18400 5800
rect 18800 -200 18900 5800
rect 17700 -300 18900 -200
rect 1900 -800 5100 -400
rect 11600 -600 11800 -300
rect 14400 -600 14600 -300
rect 11600 -800 14600 -600
<< viali >>
rect -2200 36400 -1800 42400
rect 1200 36400 1600 42400
rect -2200 29200 -1800 35200
rect 1200 29200 1600 35200
rect 2000 29200 2200 35200
rect 5400 36400 5800 42400
rect 7600 36400 9000 42400
rect 10800 36400 11200 42400
rect 6700 35700 9900 35900
rect 5400 29200 5800 35200
rect 7600 29200 7800 35200
rect 8800 29200 9000 35200
rect 10800 29200 11200 35200
rect 12900 35500 13300 36100
rect 15000 36400 15400 42400
rect 18400 36400 18800 42400
rect 14400 29200 14600 35200
rect 15000 29200 15400 35200
rect 18400 29200 18800 35200
rect 2800 21700 3000 27700
rect 6700 28500 8500 28700
rect 4800 25400 5000 27700
rect 6200 21700 6400 24200
rect 8200 21700 8400 27700
rect 10200 21700 10400 24200
rect 11600 25400 11800 27700
rect 13600 21700 13800 27700
rect 6100 21000 7300 21200
rect 2800 14500 3000 20500
rect 4800 14500 5000 16800
rect 3900 14000 4500 14200
rect 6200 18000 6400 20500
rect 8200 14500 8400 20500
rect 10200 18000 10400 20500
rect 11600 14500 11800 16800
rect 13600 14500 13800 20500
rect 12100 14000 12700 14200
rect -2200 7000 -1800 13000
rect 1200 7000 1600 13000
rect 2000 7000 2200 13000
rect -2200 -200 -1800 5800
rect 1200 -200 1600 5800
rect 3300 6100 3700 6700
rect 5400 7000 5800 13000
rect 7600 7000 7800 13000
rect 8800 7000 9000 13000
rect 10800 7000 11200 13000
rect 6700 6300 9900 6500
rect 5400 -200 5800 5800
rect 7600 -200 9000 5800
rect 10800 -200 11200 5800
rect 14400 7000 14600 13000
rect 15000 7000 15400 13000
rect 18400 7000 18800 13000
rect 15000 -200 15400 5800
rect 18400 -200 18800 5800
<< metal1 >>
rect -2500 42500 19100 42900
rect -2300 42400 -1700 42500
rect -2300 36400 -2200 42400
rect -1800 36400 -1700 42400
rect -2300 35200 -1700 36400
rect -2300 29200 -2200 35200
rect -1800 29200 -1700 35200
rect -2300 29100 -1700 29200
rect 1100 42400 1700 42500
rect 1100 36400 1200 42400
rect 1600 36400 1700 42400
rect 1100 35200 1700 36400
rect 5300 42400 5900 42500
rect 5300 36400 5400 42400
rect 5800 36400 5900 42400
rect 1100 29200 1200 35200
rect 1600 29200 1700 35200
rect 1100 29100 1700 29200
rect 1900 35200 2300 35300
rect 1900 29200 2000 35200
rect 2200 29200 2300 35200
rect 1900 29100 2300 29200
rect 5300 35200 5900 36400
rect 7500 42400 9100 42500
rect 7500 36400 7600 42400
rect 9000 36400 9100 42400
rect 7500 36300 9100 36400
rect 10700 42400 11300 42500
rect 10700 36400 10800 42400
rect 11200 36400 11300 42400
rect 6600 35900 10000 36000
rect 6600 35700 6700 35900
rect 9900 35700 10000 35900
rect 6600 35600 10000 35700
rect 5300 29200 5400 35200
rect 5800 29200 5900 35200
rect 5300 29100 5900 29200
rect 7500 35200 7900 35300
rect 7500 29200 7600 35200
rect 7800 29200 7900 35200
rect 7500 29100 7900 29200
rect 8700 35200 9100 35300
rect 8700 29200 8800 35200
rect 9000 29200 9100 35200
rect 8700 29100 9100 29200
rect 10700 35200 11300 36400
rect 14900 42400 15500 42500
rect 14900 36400 15000 42400
rect 15400 36400 15500 42400
rect 12800 36100 13400 36200
rect 12800 35500 12900 36100
rect 13300 35500 13400 36100
rect 12800 35400 13400 35500
rect 10700 29200 10800 35200
rect 11200 29200 11300 35200
rect 10700 29100 11300 29200
rect 11500 29100 11900 35300
rect 14300 35200 14700 35300
rect 14300 29200 14400 35200
rect 14600 29200 14700 35200
rect 14300 29100 14700 29200
rect 14900 35200 15500 36400
rect 14900 29200 15000 35200
rect 15400 29200 15500 35200
rect 14900 29100 15500 29200
rect 18300 42400 18900 42500
rect 18300 36400 18400 42400
rect 18800 36400 18900 42400
rect 18300 35200 18900 36400
rect 18300 29200 18400 35200
rect 18800 29200 18900 35200
rect 18300 29100 18900 29200
rect 6600 28700 8600 28800
rect 6600 28500 6700 28700
rect 8500 28500 8600 28700
rect 6600 28400 8600 28500
rect 2700 27700 3100 27800
rect 2700 21700 2800 27700
rect 3000 21700 3100 27700
rect 4700 27700 5100 27800
rect 4700 25400 4800 27700
rect 5000 25400 5100 27700
rect 4700 25300 5100 25400
rect 7500 27700 9100 27800
rect 2700 20500 3100 21700
rect 6100 24200 6500 24300
rect 6100 21700 6200 24200
rect 6400 21700 6500 24200
rect 6100 21600 6500 21700
rect 7500 21700 8200 27700
rect 8400 21700 9100 27700
rect 11500 27700 11900 27800
rect 11500 25400 11600 27700
rect 11800 25400 11900 27700
rect 11500 25300 11900 25400
rect 13500 27700 13900 27800
rect 7500 21600 9100 21700
rect 10100 24200 10500 24300
rect 10100 21700 10200 24200
rect 10400 21700 10500 24200
rect 10100 21600 10500 21700
rect 13500 21700 13600 27700
rect 13800 21700 13900 27700
rect 6000 21200 7400 21300
rect 6000 21000 6100 21200
rect 7300 21000 7400 21200
rect 6000 20900 7400 21000
rect 8100 20600 8500 21600
rect 2700 14500 2800 20500
rect 3000 14500 3100 20500
rect 6100 20500 6500 20600
rect 6100 18000 6200 20500
rect 6400 18000 6500 20500
rect 6100 17900 6500 18000
rect 7500 20500 9100 20600
rect 2700 14300 3100 14500
rect 4700 16800 5100 16900
rect 4700 14500 4800 16800
rect 5000 14500 5100 16800
rect 4700 14400 5100 14500
rect 7500 14500 8200 20500
rect 8400 14500 9100 20500
rect 10100 20500 10500 20600
rect 10100 18000 10200 20500
rect 10400 18000 10500 20500
rect 10100 17900 10500 18000
rect 13500 20500 13900 21700
rect 7500 14400 9100 14500
rect 11500 16800 11900 16900
rect 11500 14500 11600 16800
rect 11800 14500 11900 16800
rect 11500 14400 11900 14500
rect 13500 14500 13600 20500
rect 13800 14500 13900 20500
rect 8100 14300 8500 14400
rect 13500 14300 13900 14500
rect -2500 14200 19100 14300
rect -2500 14000 3900 14200
rect 4500 14000 12100 14200
rect 12700 14000 19100 14200
rect -2500 13900 19100 14000
rect -2300 13000 -1700 13100
rect -2300 7000 -2200 13000
rect -1800 7000 -1700 13000
rect -2300 5800 -1700 7000
rect -2300 -200 -2200 5800
rect -1800 -200 -1700 5800
rect -2300 -300 -1700 -200
rect 1100 13000 1700 13100
rect 1100 7000 1200 13000
rect 1600 7000 1700 13000
rect 1100 5800 1700 7000
rect 1900 13000 2300 13100
rect 1900 7000 2000 13000
rect 2200 7000 2300 13000
rect 1900 6900 2300 7000
rect 4700 6900 5100 13100
rect 5300 13000 5900 13100
rect 5300 7000 5400 13000
rect 5800 7000 5900 13000
rect 3200 6700 3800 6800
rect 3200 6100 3300 6700
rect 3700 6100 3800 6700
rect 3200 6000 3800 6100
rect 1100 -200 1200 5800
rect 1600 -200 1700 5800
rect 1100 -300 1700 -200
rect 5300 5800 5900 7000
rect 7500 13000 7900 13100
rect 7500 7000 7600 13000
rect 7800 7000 7900 13000
rect 7500 6900 7900 7000
rect 8700 13000 9100 13100
rect 8700 7000 8800 13000
rect 9000 7000 9100 13000
rect 8700 6900 9100 7000
rect 10700 13000 11300 13100
rect 10700 7000 10800 13000
rect 11200 7000 11300 13000
rect 6600 6500 10000 6600
rect 6600 6300 6700 6500
rect 9900 6300 10000 6500
rect 6600 6200 10000 6300
rect 5300 -200 5400 5800
rect 5800 -200 5900 5800
rect 5300 -300 5900 -200
rect 7500 5800 9100 5900
rect 7500 -200 7600 5800
rect 9000 -200 9100 5800
rect 7500 -300 9100 -200
rect 10700 5800 11300 7000
rect 14300 13000 14700 13100
rect 14300 7000 14400 13000
rect 14600 7000 14700 13000
rect 14300 6900 14700 7000
rect 14900 13000 15500 13100
rect 14900 7000 15000 13000
rect 15400 7000 15500 13000
rect 10700 -200 10800 5800
rect 11200 -200 11300 5800
rect 10700 -300 11300 -200
rect 14900 5800 15500 7000
rect 14900 -200 15000 5800
rect 15400 -200 15500 5800
rect 14900 -300 15500 -200
rect 18300 13000 18900 13100
rect 18300 7000 18400 13000
rect 18800 7000 18900 13000
rect 18300 5800 18900 7000
rect 18300 -200 18400 5800
rect 18800 -200 18900 5800
rect 18300 -300 18900 -200
rect -2500 -700 19100 -300
<< via1 >>
rect 2000 29200 2200 35200
rect 6700 35700 9900 35900
rect 7600 29200 7800 35200
rect 12900 35500 13300 36100
rect 14400 29200 14600 35200
rect 6700 28500 8500 28700
rect 4800 25400 5000 27700
rect 6200 21700 6400 24200
rect 11600 25400 11800 27700
rect 10200 21700 10400 24200
rect 6100 21000 7300 21200
rect 6200 18000 6400 20500
rect 4800 14500 5000 16800
rect 10200 18000 10400 20500
rect 11600 14500 11800 16800
rect 2000 7000 2200 13000
rect 3300 6100 3700 6700
rect 7600 7000 7800 13000
rect 8800 7000 9000 13000
rect 6700 6300 9900 6500
rect 14400 7000 14600 13000
<< metal2 >>
rect 12800 36100 13400 36200
rect 12800 36000 12900 36100
rect 6600 35900 12900 36000
rect 6600 35700 6700 35900
rect 9900 35700 12900 35900
rect 6600 35600 12900 35700
rect 12800 35500 12900 35600
rect 13300 35500 13400 36100
rect 12800 35400 13400 35500
rect 1900 35200 2300 35300
rect 1900 29200 2000 35200
rect 2200 29200 2300 35200
rect 1900 29100 2300 29200
rect 7500 35200 7900 35300
rect 7500 29200 7600 35200
rect 7800 29500 7900 35200
rect 14300 35200 14700 35300
rect 7800 29200 9100 29500
rect 7500 29100 9100 29200
rect 14300 29200 14400 35200
rect 14600 29200 14700 35200
rect 14300 29100 14700 29200
rect 6600 28700 8600 28800
rect 6600 28500 6700 28700
rect 8500 28500 8600 28700
rect 6600 28400 8600 28500
rect 4700 27700 5100 27800
rect 4700 25400 4800 27700
rect 5000 25400 5100 27700
rect 4700 25300 5100 25400
rect 7500 25200 7900 28400
rect -2500 24400 7900 25200
rect 6100 24200 6500 24300
rect 6100 21700 6200 24200
rect 6400 21700 6500 24200
rect -2500 21300 -1700 21700
rect 6100 21600 6500 21700
rect -2500 21200 7400 21300
rect -2500 21000 6100 21200
rect 7300 21000 7400 21200
rect -2500 20900 7400 21000
rect 6100 20500 6500 20600
rect 6100 18000 6200 20500
rect 6400 18000 6500 20500
rect 6100 17900 6500 18000
rect 4700 16800 5100 16900
rect 4700 14500 4800 16800
rect 5000 14500 5100 16800
rect 4700 14400 5100 14500
rect 1900 13000 2300 13100
rect 1900 7000 2000 13000
rect 2200 7000 2300 13000
rect 1900 6900 2300 7000
rect 7500 13000 7900 24400
rect 7500 7000 7600 13000
rect 7800 7000 7900 13000
rect 7500 6900 7900 7000
rect 8700 25200 9100 29100
rect 11500 27700 11900 27800
rect 11500 25400 11600 27700
rect 11800 25400 11900 27700
rect 11500 25300 11900 25400
rect 8700 24400 19100 25200
rect 8700 17800 9100 24400
rect 10100 24200 10500 24300
rect 10100 21700 10200 24200
rect 10400 21700 10500 24200
rect 10100 21600 10500 21700
rect 10100 20500 10500 20600
rect 10100 18000 10200 20500
rect 10400 18000 10500 20500
rect 10100 17900 10500 18000
rect 8700 17000 19100 17800
rect 8700 13000 9100 17000
rect 11500 16800 11900 16900
rect 11500 14500 11600 16800
rect 11800 14500 11900 16800
rect 11500 14400 11900 14500
rect 8700 7000 8800 13000
rect 9000 7000 9100 13000
rect 8700 6900 9100 7000
rect 14300 13000 14700 13100
rect 14300 7000 14400 13000
rect 14600 7000 14700 13000
rect 14300 6900 14700 7000
rect 3200 6700 3800 6800
rect 3200 6100 3300 6700
rect 3700 6600 3800 6700
rect 3700 6500 10000 6600
rect 3700 6300 6700 6500
rect 9900 6300 10000 6500
rect 3700 6200 10000 6300
rect 3700 6100 3800 6200
rect 3200 6000 3800 6100
<< via2 >>
rect 2000 29200 2200 35200
rect 14400 29200 14600 35200
rect 4800 25400 5000 27700
rect 6200 21700 6400 24200
rect 6200 18000 6400 20500
rect 4800 14500 5000 16800
rect 2000 7000 2200 13000
rect 11600 25400 11800 27700
rect 10200 21700 10400 24200
rect 10200 18000 10400 20500
rect 11600 14500 11800 16800
rect 14400 7000 14600 13000
<< metal3 >>
rect 1900 35200 2300 35300
rect 1900 29500 2000 35200
rect 1300 29200 2000 29500
rect 2200 29200 2300 35200
rect 1300 29100 2300 29200
rect 14300 35200 14700 35300
rect 14300 29200 14400 35200
rect 14600 29200 14700 35200
rect 1300 6700 1700 29100
rect 4700 27700 5100 27800
rect 4700 25700 4800 27700
rect 4200 25400 4800 25700
rect 5000 25400 5100 27700
rect 11500 27700 11900 27800
rect 11500 25700 11600 27700
rect 4200 25300 5100 25400
rect 11000 25400 11600 25700
rect 11800 25400 11900 27700
rect 11000 25300 11900 25400
rect 4200 14300 4600 25300
rect 6100 24200 6500 24300
rect 6100 22000 6200 24200
rect 5600 21700 6200 22000
rect 6400 21700 6500 24200
rect 10100 24200 10500 24300
rect 10100 22000 10200 24200
rect 5600 21600 6500 21700
rect 8100 21700 10200 22000
rect 10400 21700 10500 24200
rect 8100 21600 10500 21700
rect 5600 17800 6000 21600
rect 8100 20600 8500 21600
rect 6100 20500 8500 20600
rect 6100 18000 6200 20500
rect 6400 20200 8500 20500
rect 10100 20500 10500 20600
rect 6400 18000 6500 20200
rect 6100 17900 6500 18000
rect 10100 18000 10200 20500
rect 10400 18000 10500 20500
rect 10100 17800 10500 18000
rect 5600 17400 10500 17800
rect 11000 16900 11400 25300
rect 4700 16800 11400 16900
rect 4700 14500 4800 16800
rect 5000 16500 11400 16800
rect 11500 16800 11900 16900
rect 5000 14500 5100 16500
rect 4700 14400 5100 14500
rect 11500 14500 11600 16800
rect 11800 14500 11900 16800
rect 11500 14300 11900 14500
rect 4200 13900 11900 14300
rect 12000 13900 12800 14300
rect 14300 13700 14700 29200
rect 1900 13300 14700 13700
rect 1900 13000 2300 13300
rect 1900 7000 2000 13000
rect 2200 7000 2300 13000
rect 1900 6900 2300 7000
rect 14300 13000 14700 13100
rect 14300 7000 14400 13000
rect 14600 7000 14700 13000
rect 14300 6700 14700 7000
rect 1300 6300 14700 6700
<< labels >>
flabel metal2 -2500 24800 -2500 24800 0 FreeSans 1600 0 0 0 I_IN
port 0 nsew
flabel metal2 -2500 21300 -2500 21300 0 FreeSans 1600 0 0 0 VBP
port 1 nsew
flabel metal2 19100 24800 19100 24800 0 FreeSans 1600 0 0 0 I_OUT
port 2 nsew
flabel metal1 -2500 14100 -2500 14100 0 FreeSans 1600 0 0 0 VP
port 3 nsew
flabel metal1 -2500 -500 -2500 -500 0 FreeSans 1600 0 0 0 VN
port 5 nsew
<< end >>
