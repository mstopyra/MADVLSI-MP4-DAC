magic
tech sky130A
timestamp 1701150204
<< nmos >>
rect 2600 14500 3000 17700
rect 18100 14500 18500 17700
rect 19600 14500 20000 17700
rect 2600 10900 3000 14100
rect 18300 10800 18700 14000
<< ndiff >>
rect 2300 17500 2600 17700
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 2300 14500 2600 14700
rect 3000 17500 3300 17700
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14500 3300 14700
rect 17800 17500 18100 17700
rect 17800 14700 17900 17500
rect 18000 14700 18100 17500
rect 17800 14500 18100 14700
rect 18500 17500 18800 17700
rect 18500 14700 18600 17500
rect 18700 14700 18800 17500
rect 18500 14500 18800 14700
rect 19300 17500 19600 17700
rect 19300 14700 19400 17500
rect 19500 14700 19600 17500
rect 19300 14500 19600 14700
rect 20000 17500 20300 17700
rect 20000 14700 20100 17500
rect 20200 14700 20300 17500
rect 20000 14500 20300 14700
rect 2300 13900 2600 14100
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 2300 10900 2600 11100
rect 3000 13900 3300 14100
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 10900 3300 11100
rect 18000 13800 18300 14000
rect 18000 11000 18100 13800
rect 18200 11000 18300 13800
rect 18000 10800 18300 11000
rect 18700 13800 19000 14000
rect 18700 11000 18800 13800
rect 18900 11000 19000 13800
rect 18700 10800 19000 11000
<< ndiffc >>
rect 2400 14700 2500 17500
rect 3100 14700 3200 17500
rect 17900 14700 18000 17500
rect 18600 14700 18700 17500
rect 19400 14700 19500 17500
rect 20100 14700 20200 17500
rect 2400 11100 2500 13900
rect 3100 11100 3200 13900
rect 18100 11000 18200 13800
rect 18800 11000 18900 13800
<< psubdiff >>
rect 2000 17500 2300 17700
rect 2000 16210 2100 17500
rect 2002 15948 2100 16210
rect 2000 14700 2100 15948
rect 2200 14700 2300 17500
rect 2000 14500 2300 14700
rect 17530 17600 17800 17700
rect 17530 14600 17600 17600
rect 17700 14600 17800 17600
rect 17530 14500 17800 14600
rect 19000 17500 19300 17700
rect 19000 14700 19100 17500
rect 19200 14700 19300 17500
rect 19000 14500 19300 14700
rect 2000 13900 2300 14100
rect 2000 11100 2100 13900
rect 2200 11100 2300 13900
rect 2000 10900 2300 11100
rect 17700 13800 18000 14000
rect 17700 11000 17800 13800
rect 17900 11000 18000 13800
rect 17700 10800 18000 11000
<< psubdiffcont >>
rect 2100 14700 2200 17500
rect 17600 14600 17700 17600
rect 19100 14700 19200 17500
rect 2100 11100 2200 13900
rect 17800 11000 17900 13800
<< poly >>
rect 2600 17700 3000 18000
rect 17200 17950 18500 18000
rect 17200 17850 18150 17950
rect 18450 17850 18500 17950
rect 17200 17800 18500 17850
rect 19200 17950 20000 18000
rect 19200 17850 19250 17950
rect 19450 17850 20000 17950
rect 19200 17800 20000 17850
rect 18100 17700 18500 17800
rect 19600 17700 20000 17800
rect 2600 14350 3000 14500
rect 18100 14400 18500 14500
rect 2600 14250 2650 14350
rect 2950 14250 3000 14350
rect 19600 14300 20000 14500
rect 2600 14100 3000 14250
rect 18300 14100 20000 14300
rect 18300 14000 18700 14100
rect 2600 10800 3000 10900
rect 18300 10700 18700 10800
<< polycont >>
rect 18150 17850 18450 17950
rect 19250 17850 19450 17950
rect 2650 14250 2950 14350
<< locali >>
rect 2000 17800 3500 18000
rect 17600 17600 17700 18000
rect 18100 17950 18500 18000
rect 18100 17850 18150 17950
rect 18450 17850 18500 17950
rect 18100 17800 18500 17850
rect 19200 17950 19500 18000
rect 19200 17850 19250 17950
rect 19450 17850 19500 17950
rect 19200 17600 19500 17850
rect 2000 17500 2600 17600
rect 2000 16210 2100 17500
rect 2002 15948 2100 16210
rect 2000 14700 2100 15948
rect 2200 14700 2400 17500
rect 2500 14700 2600 17500
rect 2000 14600 2600 14700
rect 3000 17500 3300 17600
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14600 3300 14700
rect 17800 17500 18100 17600
rect 17800 14700 17900 17500
rect 18000 14700 18100 17500
rect 17800 14600 18100 14700
rect 18500 17500 18800 17600
rect 18500 14700 18600 17500
rect 18700 14700 18800 17500
rect 18500 14600 18800 14700
rect 19000 17500 19600 17600
rect 19000 14700 19100 17500
rect 19200 14700 19400 17500
rect 19500 14700 19600 17500
rect 19000 14600 19600 14700
rect 20000 17500 20300 17600
rect 20000 14700 20100 17500
rect 20200 14700 20300 17500
rect 20000 14600 20300 14700
rect 2400 14400 2500 14600
rect 2400 14350 3000 14400
rect 2400 14250 2650 14350
rect 2950 14250 3000 14350
rect 2400 14200 3000 14250
rect 17600 14300 17700 14600
rect 18500 14500 18700 14600
rect 20000 14500 20200 14600
rect 17600 14200 17900 14300
rect 2400 14000 2500 14200
rect 2000 13900 2600 14000
rect 2000 11100 2100 13900
rect 2200 11100 2400 13900
rect 2500 11100 2600 13900
rect 2000 11000 2600 11100
rect 3000 13900 3300 14000
rect 17800 13900 17900 14200
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 11000 3300 11100
rect 17700 13800 18300 13900
rect 17700 11000 17800 13800
rect 17900 11000 18100 13800
rect 18200 11000 18300 13800
rect 17200 10900 17500 11000
rect 17700 10900 18300 11000
rect 18700 13800 19000 13900
rect 18700 11000 18800 13800
rect 18900 11000 19000 13800
rect 18700 10900 19000 11000
rect 17300 10700 17500 10900
rect 18700 10800 18900 10900
rect 17250 10650 17450 10700
rect 17250 10500 17300 10650
rect 17400 10600 17450 10650
<< viali >>
rect 2400 14700 2500 17500
rect 3100 16000 3200 16200
rect 17900 16000 18000 16200
rect 18600 15000 18700 15200
rect 19400 14700 19500 17500
rect 20100 15950 20200 16250
rect 2400 11100 2500 13900
rect 3100 12200 3200 12400
rect 18100 11000 18200 13800
rect 18800 12150 18900 12450
rect 17300 10550 17400 10650
<< metal1 >>
rect 2300 17500 2600 17600
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 19300 17500 19600 17600
rect 19300 16300 19400 17500
rect 3050 16200 3500 16300
rect 3050 16000 3100 16200
rect 3200 16000 3500 16200
rect 3050 15900 3500 16000
rect 17500 16200 18400 16300
rect 17500 16000 17900 16200
rect 18000 16000 18400 16200
rect 17500 15900 18400 16000
rect 19000 15900 19400 16300
rect 18500 15200 18800 15300
rect 18500 15000 18600 15200
rect 18700 15000 18800 15200
rect 18500 14900 18800 15000
rect 2300 13900 2600 14700
rect 19300 14700 19400 15900
rect 19500 14700 19600 17500
rect 20000 16250 20250 16300
rect 20000 15950 20100 16250
rect 20200 15950 20250 16250
rect 20000 15900 20250 15950
rect 19300 14500 19600 14700
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 18000 14100 19600 14500
rect 18000 13800 18700 14100
rect 3000 12400 3500 12500
rect 3000 12200 3100 12400
rect 3200 12200 3500 12400
rect 3000 12100 3500 12200
rect 17500 12450 17700 12500
rect 17500 12150 17550 12450
rect 17650 12150 17700 12450
rect 17500 12100 17700 12150
rect 2300 10000 2600 11100
rect 18000 11000 18100 13800
rect 18200 11000 18700 13800
rect 18750 12450 18950 12500
rect 18750 12150 18800 12450
rect 18900 12150 18950 12450
rect 18750 12100 18950 12150
rect 17250 10650 17300 10700
rect 17000 10550 17300 10650
rect 17250 10500 17300 10550
rect 18000 10000 18700 11000
rect 2300 6800 3500 10000
rect 17500 6800 18700 10000
<< via1 >>
rect 3100 16000 3200 16200
rect 17900 16000 18000 16200
rect 18600 15000 18700 15200
rect 20100 15950 20200 16250
rect 3100 12200 3200 12400
rect 17550 12150 17650 12450
rect 18800 12150 18900 12450
rect 17300 10550 17400 10650
<< metal2 >>
rect 2000 16210 3300 16300
rect 2002 16200 3300 16210
rect 2002 16000 3100 16200
rect 3200 16000 3300 16200
rect 2002 15948 3300 16000
rect 2000 15900 3300 15948
rect 17800 16250 20250 16300
rect 17800 16200 20100 16250
rect 17800 16000 17900 16200
rect 18000 16000 20100 16200
rect 17800 15950 20100 16000
rect 20200 15950 20250 16250
rect 17800 15900 20250 15950
rect 17100 15200 20900 15300
rect 17100 15000 18600 15200
rect 18700 15000 20900 15200
rect 17100 14900 20900 15000
rect 2000 12400 3300 12500
rect 2000 12200 3100 12400
rect 3200 12200 3300 12400
rect 2000 12100 3300 12200
rect 17100 10700 17400 14900
rect 17500 12450 20900 12500
rect 17500 12150 17550 12450
rect 17650 12150 18800 12450
rect 18900 12150 20900 12450
rect 17500 12100 20900 12150
rect 17250 10650 17450 10700
rect 17250 10550 17300 10650
rect 17400 10550 17450 10650
rect 17250 10500 17450 10550
use DAC_block  DAC_block_14
timestamp 1701149695
transform 1 0 1800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_15
timestamp 1701149695
transform 1 0 13800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_16
timestamp 1701149695
transform 1 0 3800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_17
timestamp 1701149695
transform 1 0 5800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_18
timestamp 1701149695
transform 1 0 7800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_19
timestamp 1701149695
transform 1 0 9800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_20
timestamp 1701149695
transform 1 0 11800 0 1 10700
box 1700 -10800 3700 7300
<< labels >>
flabel metal2 2000 12300 2000 12300 0 FreeSans 800 0 0 0 I_OUT
port 3 nsew
flabel space 4800 -100 4800 -100 0 FreeSans 800 0 0 0 D_6
port 5 nsew
flabel space 6800 -100 6800 -100 0 FreeSans 800 0 0 0 D_5
port 6 nsew
flabel space 8800 -100 8800 -100 0 FreeSans 800 0 0 0 D_4
port 7 nsew
flabel space 10800 -100 10800 -100 0 FreeSans 800 0 0 0 D_3
port 8 nsew
flabel space 12800 -100 12800 -100 0 FreeSans 800 0 0 0 D_2
port 9 nsew
flabel space 14800 -100 14800 -100 0 FreeSans 800 0 0 0 D_1
port 10 nsew
flabel space 16800 -100 16800 -100 0 FreeSans 800 0 0 0 D_0
port 11 nsew
flabel metal2 20900 12300 20900 12300 0 FreeSans 800 0 0 0 I_OUT_LD
port 14 nsew
flabel metal1 2300 8300 2300 8300 0 FreeSans 800 0 0 0 VN
port 16 nsew
flabel space 3500 3300 3500 3300 0 FreeSans 800 0 0 0 VP
port 18 nsew
flabel locali 2000 17900 2000 17900 0 FreeSans 800 0 0 0 I_IN
port 17 nsew
flabel metal2 20900 15100 20900 15100 0 FreeSans 800 0 0 0 I_DUMP
port 12 nsew
<< end >>
