magic
tech sky130A
timestamp 1701144982
<< nwell >>
rect -1250 14150 9550 21550
rect 3050 10500 3650 10600
rect -1250 -450 9550 6950
<< nmos >>
rect 1900 10750 2300 13950
rect 2600 10750 3000 13950
rect 3300 10750 3700 13950
rect 4600 10750 5000 13950
rect 5300 10750 5700 13950
rect 6000 10750 6400 13950
rect 1900 7150 2300 10350
rect 2600 7150 3000 10350
rect 3300 7150 3700 10350
rect 4600 7150 5000 10350
rect 5300 7150 5700 10350
rect 6000 7150 6400 10350
<< pmos >>
rect -500 18100 -100 21300
rect 1200 18100 1600 21300
rect 1900 18100 2300 21300
rect 3300 18100 3700 21300
rect 4600 18100 5000 21300
rect 6000 18100 6400 21300
rect 6700 18100 7100 21300
rect 8400 18100 8800 21300
rect -500 14500 -100 17700
rect 1200 14500 1600 17700
rect 1900 14500 2300 17700
rect 3300 14500 3700 17700
rect 4600 14500 5000 17700
rect 6000 14500 6400 17700
rect 6700 14500 7100 17700
rect 8400 14500 8800 17700
rect -500 3400 -100 6600
rect 1200 3400 1600 6600
rect 1900 3400 2300 6600
rect 3300 3400 3700 6600
rect 4600 3400 5000 6600
rect 6000 3400 6400 6600
rect 6700 3400 7100 6600
rect 8400 3400 8800 6600
rect -500 -200 -100 3000
rect 1200 -200 1600 3000
rect 1900 -200 2300 3000
rect 3300 -200 3700 3000
rect 4600 -200 5000 3000
rect 6000 -200 6400 3000
rect 6700 -200 7100 3000
rect 8400 -200 8800 3000
<< ndiff >>
rect 1600 13850 1900 13950
rect 1600 10850 1700 13850
rect 1800 10850 1900 13850
rect 1600 10750 1900 10850
rect 2300 13850 2600 13950
rect 2300 10850 2400 13850
rect 2500 10850 2600 13850
rect 2300 10750 2600 10850
rect 3000 13850 3300 13950
rect 3000 10850 3100 13850
rect 3200 10850 3300 13850
rect 3000 10750 3300 10850
rect 3700 13850 4000 13950
rect 4300 13850 4600 13950
rect 3700 10850 3800 13850
rect 3900 10850 4000 13850
rect 4300 10850 4400 13850
rect 4500 10850 4600 13850
rect 3700 10750 4000 10850
rect 4300 10750 4600 10850
rect 5000 13800 5300 13950
rect 5000 10850 5100 13800
rect 5200 10850 5300 13800
rect 5000 10750 5300 10850
rect 5700 13850 6000 13950
rect 5700 10850 5800 13850
rect 5900 10850 6000 13850
rect 5700 10750 6000 10850
rect 6400 13850 6700 13950
rect 6400 10850 6500 13850
rect 6600 10850 6700 13850
rect 6400 10750 6700 10850
rect 1600 10250 1900 10350
rect 1600 7250 1700 10250
rect 1800 7250 1900 10250
rect 1600 7150 1900 7250
rect 2300 10250 2600 10350
rect 2300 7250 2400 10250
rect 2500 7250 2600 10250
rect 2300 7150 2600 7250
rect 3000 10250 3300 10350
rect 3000 7250 3100 10250
rect 3200 7250 3300 10250
rect 3000 7150 3300 7250
rect 3700 10250 4000 10350
rect 4300 10250 4600 10350
rect 3700 7250 3800 10250
rect 3900 7250 4000 10250
rect 4300 7250 4400 10250
rect 4500 7250 4600 10250
rect 3700 7150 4000 7250
rect 4300 7150 4600 7250
rect 5000 10250 5300 10350
rect 5000 7250 5100 10250
rect 5200 7250 5300 10250
rect 5000 7150 5300 7250
rect 5700 10250 6000 10350
rect 5700 7250 5800 10250
rect 5900 7250 6000 10250
rect 5700 7150 6000 7250
rect 6400 10250 6700 10350
rect 6400 7250 6500 10250
rect 6600 7250 6700 10250
rect 6400 7150 6700 7250
<< pdiff >>
rect -800 21200 -500 21300
rect -800 18200 -700 21200
rect -600 18200 -500 21200
rect -800 18100 -500 18200
rect -100 21200 200 21300
rect -100 18200 0 21200
rect 100 18200 200 21200
rect -100 18100 200 18200
rect 900 21200 1200 21300
rect 900 18200 1000 21200
rect 1100 18200 1200 21200
rect 900 18100 1200 18200
rect 1600 21200 1900 21300
rect 1600 18200 1700 21200
rect 1800 18200 1900 21200
rect 1600 18100 1900 18200
rect 2300 21200 2600 21300
rect 3000 21200 3300 21300
rect 2300 18200 2400 21200
rect 2500 18200 2600 21200
rect 3000 18200 3100 21200
rect 3200 18200 3300 21200
rect 2300 18100 2600 18200
rect 3000 18100 3300 18200
rect 3700 21200 4600 21300
rect 3700 18200 3800 21200
rect 4500 18200 4600 21200
rect 3700 18100 4600 18200
rect 5000 21200 5300 21300
rect 5700 21200 6000 21300
rect 5000 18200 5100 21200
rect 5200 18200 5300 21200
rect 5700 18200 5800 21200
rect 5900 18200 6000 21200
rect 5000 18100 5300 18200
rect 5700 18100 6000 18200
rect 6400 21200 6700 21300
rect 6400 18200 6500 21200
rect 6600 18200 6700 21200
rect 6400 18100 6700 18200
rect 7100 21200 7400 21300
rect 7100 18200 7200 21200
rect 7300 18200 7400 21200
rect 7100 18100 7400 18200
rect 8100 21200 8400 21300
rect 8100 18200 8200 21200
rect 8300 18200 8400 21200
rect 8100 18100 8400 18200
rect 8800 21200 9100 21300
rect 8800 18200 8900 21200
rect 9000 18200 9100 21200
rect 8800 18100 9100 18200
rect -800 17600 -500 17700
rect -800 14600 -700 17600
rect -600 14600 -500 17600
rect -800 14500 -500 14600
rect -100 17600 200 17700
rect -100 14600 0 17600
rect 100 14600 200 17600
rect -100 14500 200 14600
rect 900 17600 1200 17700
rect 900 14600 1000 17600
rect 1100 14600 1200 17600
rect 900 14500 1200 14600
rect 1600 17600 1900 17700
rect 1600 14600 1700 17600
rect 1800 14600 1900 17600
rect 1600 14500 1900 14600
rect 2300 17600 2600 17700
rect 3000 17600 3300 17700
rect 2300 14600 2400 17600
rect 2500 14600 2600 17600
rect 3000 14600 3100 17600
rect 3200 14600 3300 17600
rect 2300 14500 2600 14600
rect 3000 14500 3300 14600
rect 3700 17600 4000 17700
rect 3700 14600 3800 17600
rect 3900 14600 4000 17600
rect 3700 14500 4000 14600
rect 4300 17600 4600 17700
rect 4300 14600 4400 17600
rect 4500 14600 4600 17600
rect 4300 14500 4600 14600
rect 5000 17600 5300 17700
rect 5700 17600 6000 17700
rect 5000 14600 5100 17600
rect 5200 14600 5300 17600
rect 5700 14600 5800 17600
rect 5900 14600 6000 17600
rect 5000 14500 5300 14600
rect 5700 14500 6000 14600
rect 6400 17600 6700 17700
rect 6400 14600 6500 17600
rect 6600 14600 6700 17600
rect 6400 14500 6700 14600
rect 7100 17600 7400 17700
rect 7100 14600 7200 17600
rect 7300 14600 7400 17600
rect 7100 14500 7400 14600
rect 8100 17600 8400 17700
rect 8100 14600 8200 17600
rect 8300 14600 8400 17600
rect 8100 14500 8400 14600
rect 8800 17600 9100 17700
rect 8800 14600 8900 17600
rect 9000 14600 9100 17600
rect 8800 14500 9100 14600
rect -800 6500 -500 6600
rect -800 3500 -700 6500
rect -600 3500 -500 6500
rect -800 3400 -500 3500
rect -100 6500 200 6600
rect -100 3500 0 6500
rect 100 3500 200 6500
rect -100 3400 200 3500
rect 900 6500 1200 6600
rect 900 3500 1000 6500
rect 1100 3500 1200 6500
rect 900 3400 1200 3500
rect 1600 6500 1900 6600
rect 1600 3500 1700 6500
rect 1800 3500 1900 6500
rect 1600 3400 1900 3500
rect 2300 6500 2600 6600
rect 3000 6500 3300 6600
rect 2300 3500 2400 6500
rect 2500 3500 2600 6500
rect 3000 3500 3100 6500
rect 3200 3500 3300 6500
rect 2300 3400 2600 3500
rect 3000 3400 3300 3500
rect 3700 6500 4000 6600
rect 3700 3500 3800 6500
rect 3900 3500 4000 6500
rect 3700 3400 4000 3500
rect 4300 6500 4600 6600
rect 4300 3500 4400 6500
rect 4500 3500 4600 6500
rect 4300 3400 4600 3500
rect 5000 6500 5300 6600
rect 5700 6500 6000 6600
rect 5000 3500 5100 6500
rect 5200 3500 5300 6500
rect 5700 3500 5800 6500
rect 5900 3500 6000 6500
rect 5000 3400 5300 3500
rect 5700 3400 6000 3500
rect 6400 6500 6700 6600
rect 6400 3500 6500 6500
rect 6600 3500 6700 6500
rect 6400 3400 6700 3500
rect 7100 6500 7400 6600
rect 7100 3500 7200 6500
rect 7300 3500 7400 6500
rect 7100 3400 7400 3500
rect 8100 6500 8400 6600
rect 8100 3500 8200 6500
rect 8300 3500 8400 6500
rect 8100 3400 8400 3500
rect 8800 6500 9100 6600
rect 8800 3500 8900 6500
rect 9000 3500 9100 6500
rect 8800 3400 9100 3500
rect -800 2900 -500 3000
rect -800 -100 -700 2900
rect -600 -100 -500 2900
rect -800 -200 -500 -100
rect -100 2900 200 3000
rect -100 -100 0 2900
rect 100 -100 200 2900
rect -100 -200 200 -100
rect 900 2900 1200 3000
rect 900 -100 1000 2900
rect 1100 -100 1200 2900
rect 900 -200 1200 -100
rect 1600 2900 1900 3000
rect 1600 -100 1700 2900
rect 1800 -100 1900 2900
rect 1600 -200 1900 -100
rect 2300 2900 2600 3000
rect 3000 2900 3300 3000
rect 2300 -100 2400 2900
rect 2500 -100 2600 2900
rect 3000 -100 3100 2900
rect 3200 -100 3300 2900
rect 2300 -200 2600 -100
rect 3000 -200 3300 -100
rect 3700 2900 4600 3000
rect 3700 -100 3800 2900
rect 4500 -100 4600 2900
rect 3700 -200 4600 -100
rect 5000 2900 5300 3000
rect 5700 2900 6000 3000
rect 5000 -100 5100 2900
rect 5200 -100 5300 2900
rect 5700 -100 5800 2900
rect 5900 -100 6000 2900
rect 5000 -200 5300 -100
rect 5700 -200 6000 -100
rect 6400 2900 6700 3000
rect 6400 -100 6500 2900
rect 6600 -100 6700 2900
rect 6400 -200 6700 -100
rect 7100 2900 7400 3000
rect 7100 -100 7200 2900
rect 7300 -100 7400 2900
rect 7100 -200 7400 -100
rect 8100 2900 8400 3000
rect 8100 -100 8200 2900
rect 8300 -100 8400 2900
rect 8100 -200 8400 -100
rect 8800 2900 9100 3000
rect 8800 -100 8900 2900
rect 9000 -100 9100 2900
rect 8800 -200 9100 -100
<< ndiffc >>
rect 1700 10850 1800 13850
rect 2400 10850 2500 13850
rect 3100 10850 3200 13850
rect 3800 10850 3900 13850
rect 4400 10850 4500 13850
rect 5100 10850 5200 13800
rect 5800 10850 5900 13850
rect 6500 10850 6600 13850
rect 1700 7250 1800 10250
rect 2400 7250 2500 10250
rect 3100 7250 3200 10250
rect 3800 7250 3900 10250
rect 4400 7250 4500 10250
rect 5100 7250 5200 10250
rect 5800 7250 5900 10250
rect 6500 7250 6600 10250
<< pdiffc >>
rect -700 18200 -600 21200
rect 0 18200 100 21200
rect 1000 18200 1100 21200
rect 1700 18200 1800 21200
rect 2400 18200 2500 21200
rect 3100 18200 3200 21200
rect 3800 18200 4500 21200
rect 5100 18200 5200 21200
rect 5800 18200 5900 21200
rect 6500 18200 6600 21200
rect 7200 18200 7300 21200
rect 8200 18200 8300 21200
rect 8900 18200 9000 21200
rect -700 14600 -600 17600
rect 0 14600 100 17600
rect 1000 14600 1100 17600
rect 1700 14600 1800 17600
rect 2400 14600 2500 17600
rect 3100 14600 3200 17600
rect 3800 14600 3900 17600
rect 4400 14600 4500 17600
rect 5100 14600 5200 17600
rect 5800 14600 5900 17600
rect 6500 14600 6600 17600
rect 7200 14600 7300 17600
rect 8200 14600 8300 17600
rect 8900 14600 9000 17600
rect -700 3500 -600 6500
rect 0 3500 100 6500
rect 1000 3500 1100 6500
rect 1700 3500 1800 6500
rect 2400 3500 2500 6500
rect 3100 3500 3200 6500
rect 3800 3500 3900 6500
rect 4400 3500 4500 6500
rect 5100 3500 5200 6500
rect 5800 3500 5900 6500
rect 6500 3500 6600 6500
rect 7200 3500 7300 6500
rect 8200 3500 8300 6500
rect 8900 3500 9000 6500
rect -700 -100 -600 2900
rect 0 -100 100 2900
rect 1000 -100 1100 2900
rect 1700 -100 1800 2900
rect 2400 -100 2500 2900
rect 3100 -100 3200 2900
rect 3800 -100 4500 2900
rect 5100 -100 5200 2900
rect 5800 -100 5900 2900
rect 6500 -100 6600 2900
rect 7200 -100 7300 2900
rect 8200 -100 8300 2900
rect 8900 -100 9000 2900
<< psubdiff >>
rect 1300 13850 1600 13950
rect 1300 10850 1400 13850
rect 1500 10850 1600 13850
rect 1300 10750 1600 10850
rect 4000 13850 4300 13950
rect 4000 10850 4100 13850
rect 4200 10850 4300 13850
rect 4000 10750 4300 10850
rect 6700 13850 7000 13950
rect 6700 10850 6800 13850
rect 6900 10850 7000 13850
rect 6700 10750 7000 10850
rect 1300 10250 1600 10350
rect 1300 7250 1400 10250
rect 1500 7250 1600 10250
rect 1300 7150 1600 7250
rect 4000 10250 4300 10350
rect 4000 7250 4100 10250
rect 4200 7250 4300 10250
rect 4000 7150 4300 7250
rect 6700 10250 7000 10350
rect 6700 7250 6800 10250
rect 6900 7250 7000 10250
rect 6700 7150 7000 7250
<< nsubdiff >>
rect -1200 21200 -800 21300
rect -1200 18200 -1100 21200
rect -900 18200 -800 21200
rect -1200 18100 -800 18200
rect 500 21200 900 21300
rect 500 18200 600 21200
rect 800 18200 900 21200
rect 500 18100 900 18200
rect 2600 21200 3000 21300
rect 2600 18200 2700 21200
rect 2900 18200 3000 21200
rect 2600 18100 3000 18200
rect 5300 21200 5700 21300
rect 5300 18200 5400 21200
rect 5600 18200 5700 21200
rect 5300 18100 5700 18200
rect 7400 21200 7800 21300
rect 7400 18200 7500 21200
rect 7700 18200 7800 21200
rect 7400 18100 7800 18200
rect 9100 21200 9500 21300
rect 9100 18200 9200 21200
rect 9400 18200 9500 21200
rect 9100 18100 9500 18200
rect -1200 17600 -800 17700
rect -1200 14600 -1100 17600
rect -900 14600 -800 17600
rect -1200 14500 -800 14600
rect 500 17600 900 17700
rect 500 14600 600 17600
rect 800 14600 900 17600
rect 500 14500 900 14600
rect 2600 17600 3000 17700
rect 2600 14600 2700 17600
rect 2900 14600 3000 17600
rect 2600 14500 3000 14600
rect 5300 17600 5700 17700
rect 5300 14600 5400 17600
rect 5600 14600 5700 17600
rect 5300 14500 5700 14600
rect 7400 17600 7800 17700
rect 7400 14600 7500 17600
rect 7700 14600 7800 17600
rect 7400 14500 7800 14600
rect 9100 17600 9500 17700
rect 9100 14600 9200 17600
rect 9400 14600 9500 17600
rect 9100 14500 9500 14600
rect -1200 6500 -800 6600
rect -1200 3500 -1100 6500
rect -900 3500 -800 6500
rect -1200 3400 -800 3500
rect 500 6500 900 6600
rect 500 3500 600 6500
rect 800 3500 900 6500
rect 500 3400 900 3500
rect 2600 6500 3000 6600
rect 2600 3500 2700 6500
rect 2900 3500 3000 6500
rect 2600 3400 3000 3500
rect 5300 6500 5700 6600
rect 5300 3500 5400 6500
rect 5600 3500 5700 6500
rect 5300 3400 5700 3500
rect 7400 6500 7800 6600
rect 7400 3500 7500 6500
rect 7700 3500 7800 6500
rect 7400 3400 7800 3500
rect 9100 6500 9500 6600
rect 9100 3500 9200 6500
rect 9400 3500 9500 6500
rect 9100 3400 9500 3500
rect -1200 2900 -800 3000
rect -1200 -100 -1100 2900
rect -900 -100 -800 2900
rect -1200 -200 -800 -100
rect 500 2900 900 3000
rect 500 -100 600 2900
rect 800 -100 900 2900
rect 500 -200 900 -100
rect 2600 2900 3000 3000
rect 2600 -100 2700 2900
rect 2900 -100 3000 2900
rect 2600 -200 3000 -100
rect 5300 2900 5700 3000
rect 5300 -100 5400 2900
rect 5600 -100 5700 2900
rect 5300 -200 5700 -100
rect 7400 2900 7800 3000
rect 7400 -100 7500 2900
rect 7700 -100 7800 2900
rect 7400 -200 7800 -100
rect 9100 2900 9500 3000
rect 9100 -100 9200 2900
rect 9400 -100 9500 2900
rect 9100 -200 9500 -100
<< psubdiffcont >>
rect 1400 10850 1500 13850
rect 4100 10850 4200 13850
rect 6800 10850 6900 13850
rect 1400 7250 1500 10250
rect 4100 7250 4200 10250
rect 6800 7250 6900 10250
<< nsubdiffcont >>
rect -1100 18200 -900 21200
rect 600 18200 800 21200
rect 2700 18200 2900 21200
rect 5400 18200 5600 21200
rect 7500 18200 7700 21200
rect 9200 18200 9400 21200
rect -1100 14600 -900 17600
rect 600 14600 800 17600
rect 2700 14600 2900 17600
rect 5400 14600 5600 17600
rect 7500 14600 7700 17600
rect 9200 14600 9400 17600
rect -1100 3500 -900 6500
rect 600 3500 800 6500
rect 2700 3500 2900 6500
rect 5400 3500 5600 6500
rect 7500 3500 7700 6500
rect 9200 3500 9400 6500
rect -1100 -100 -900 2900
rect 600 -100 800 2900
rect 2700 -100 2900 2900
rect 5400 -100 5600 2900
rect 7500 -100 7700 2900
rect 9200 -100 9400 2900
<< poly >>
rect -500 21300 -100 21400
rect 1200 21300 1600 21400
rect 1900 21300 2300 21400
rect 3300 21300 3700 21400
rect 4600 21300 5000 21400
rect 6000 21300 6400 21400
rect 6700 21300 7100 21400
rect 8400 21300 8800 21400
rect -500 18050 -100 18100
rect -500 17950 -450 18050
rect -150 17950 -100 18050
rect -500 17900 -100 17950
rect -500 17700 -100 17800
rect 1200 17700 1600 18100
rect 1900 17700 2300 18100
rect 3300 18000 3700 18100
rect 4600 18000 5000 18100
rect 3300 17950 5000 18000
rect 3300 17850 3350 17950
rect 4950 17850 5000 17950
rect 3300 17800 5000 17850
rect 3300 17700 3700 17750
rect 4600 17700 5000 17750
rect 6000 17700 6400 18100
rect 6700 17700 7100 18100
rect 8400 18050 8800 18100
rect 8400 17950 8450 18050
rect 8750 17950 8800 18050
rect 8400 17900 8800 17950
rect 8400 17700 8800 17800
rect -500 14450 -100 14500
rect -500 14350 -450 14450
rect -150 14350 -100 14450
rect -500 14300 -100 14350
rect 1200 14450 1600 14500
rect 1200 14350 1250 14450
rect 1550 14350 1600 14450
rect 1200 14300 1600 14350
rect 1900 14450 2300 14500
rect 1900 14350 1950 14450
rect 2250 14350 2300 14450
rect 1900 14300 2300 14350
rect 3300 14400 3700 14500
rect 4600 14400 5000 14500
rect 3300 14350 5000 14400
rect 3300 14250 3350 14350
rect 4950 14250 5000 14350
rect 6000 14450 6400 14500
rect 6000 14350 6050 14450
rect 6350 14350 6400 14450
rect 6000 14300 6400 14350
rect 6700 14450 7100 14500
rect 6700 14350 6750 14450
rect 7050 14350 7100 14450
rect 6700 14300 7100 14350
rect 8400 14450 8800 14500
rect 8400 14350 8450 14450
rect 8750 14350 8800 14450
rect 8400 14300 8800 14350
rect 3300 14200 5000 14250
rect 1900 13950 2300 14000
rect 2600 13950 3000 14000
rect 3300 13950 3700 14000
rect 4600 13950 5000 14000
rect 5300 13950 5700 14000
rect 6000 13950 6400 14000
rect 1900 10350 2300 10750
rect 2600 10650 3000 10750
rect 3300 10650 3700 10750
rect 4600 10650 5000 10750
rect 5300 10650 5700 10750
rect 2600 10600 5700 10650
rect 2600 10500 3050 10600
rect 3650 10500 5700 10600
rect 2600 10450 5700 10500
rect 2600 10350 3000 10450
rect 3300 10350 3700 10450
rect 4600 10350 5000 10450
rect 5300 10350 5700 10450
rect 6000 10350 6400 10750
rect 1900 7100 2300 7150
rect 2600 7100 3000 7150
rect 3300 7100 3700 7150
rect 4600 7100 5000 7150
rect 5300 7100 5700 7150
rect 6000 7100 6400 7150
rect 1900 7000 1950 7100
rect 2250 7000 2300 7100
rect 1900 6950 2300 7000
rect 6000 7000 6050 7100
rect 6350 7000 6400 7100
rect 6000 6950 6400 7000
rect 3300 6850 5000 6900
rect -500 6750 -100 6800
rect -500 6650 -450 6750
rect -150 6650 -100 6750
rect -500 6600 -100 6650
rect 1200 6750 1600 6800
rect 1200 6650 1250 6750
rect 1550 6650 1600 6750
rect 1200 6600 1600 6650
rect 1900 6750 2300 6800
rect 1900 6650 1950 6750
rect 2250 6650 2300 6750
rect 1900 6600 2300 6650
rect 3300 6750 3350 6850
rect 4950 6750 5000 6850
rect 3300 6700 5000 6750
rect 3300 6600 3700 6700
rect 4600 6600 5000 6700
rect 6000 6750 6400 6800
rect 6000 6650 6050 6750
rect 6350 6650 6400 6750
rect 6000 6600 6400 6650
rect 6700 6750 7100 6800
rect 6700 6650 6750 6750
rect 7050 6650 7100 6750
rect 6700 6600 7100 6650
rect 8400 6750 8800 6800
rect 8400 6650 8450 6750
rect 8750 6650 8800 6750
rect 8400 6600 8800 6650
rect -500 3300 -100 3400
rect -500 3150 -100 3200
rect -500 3050 -450 3150
rect -150 3050 -100 3150
rect -500 3000 -100 3050
rect 1200 3000 1600 3400
rect 1900 3000 2300 3400
rect 3300 3350 3700 3400
rect 4600 3350 5000 3400
rect 3300 3250 5000 3300
rect 3300 3150 3350 3250
rect 4950 3150 5000 3250
rect 3300 3100 5000 3150
rect 3300 3000 3700 3100
rect 4600 3000 5000 3100
rect 6000 3000 6400 3400
rect 6700 3000 7100 3400
rect 8400 3300 8800 3400
rect 8400 3150 8800 3200
rect 8400 3050 8450 3150
rect 8750 3050 8800 3150
rect 8400 3000 8800 3050
rect -500 -300 -100 -200
rect 1200 -300 1600 -200
rect 1900 -300 2300 -200
rect 3300 -300 3700 -200
rect 4600 -300 5000 -200
rect 6000 -300 6400 -200
rect 6700 -300 7100 -200
rect 8400 -300 8800 -200
<< polycont >>
rect -450 17950 -150 18050
rect 3350 17850 4950 17950
rect 8450 17950 8750 18050
rect -450 14350 -150 14450
rect 1250 14350 1550 14450
rect 1950 14350 2250 14450
rect 3350 14250 4950 14350
rect 6050 14350 6350 14450
rect 6750 14350 7050 14450
rect 8450 14350 8750 14450
rect 3050 10500 3650 10600
rect 1950 7000 2250 7100
rect 6050 7000 6350 7100
rect -450 6650 -150 6750
rect 1250 6650 1550 6750
rect 1950 6650 2250 6750
rect 3350 6750 4950 6850
rect 6050 6650 6350 6750
rect 6750 6650 7050 6750
rect 8450 6650 8750 6750
rect -450 3050 -150 3150
rect 3350 3150 4950 3250
rect 8450 3050 8750 3150
<< locali >>
rect 950 21300 2550 21500
rect -1150 21200 -550 21250
rect -1150 18200 -1100 21200
rect -900 18200 -700 21200
rect -600 18200 -550 21200
rect -1150 18100 -550 18200
rect -50 21200 150 21250
rect -50 18200 0 21200
rect 100 18200 150 21200
rect -1150 18050 -100 18100
rect -1150 17950 -450 18050
rect -150 17950 -100 18050
rect -1150 17900 -100 17950
rect -50 18000 150 18200
rect 550 21200 850 21250
rect 550 18200 600 21200
rect 800 18200 850 21200
rect 550 18150 850 18200
rect 950 21200 1150 21300
rect 950 18200 1000 21200
rect 1100 18200 1150 21200
rect 950 18000 1150 18200
rect -1150 17600 -550 17900
rect -1150 14600 -1100 17600
rect -900 14600 -700 17600
rect -600 14600 -550 17600
rect -1150 14500 -550 14600
rect -50 17800 1150 18000
rect -50 17600 150 17800
rect -50 14600 0 17600
rect 100 14600 150 17600
rect -50 14500 150 14600
rect 550 17600 850 17650
rect 550 14600 600 17600
rect 800 14600 850 17600
rect 550 14550 850 14600
rect 950 17600 1150 17800
rect 950 14600 1000 17600
rect 1100 14600 1150 17600
rect 950 14550 1150 14600
rect 1650 21200 1850 21250
rect 1650 18200 1700 21200
rect 1800 18200 1850 21200
rect 1650 17600 1850 18200
rect 1650 14600 1700 17600
rect 1800 14600 1850 17600
rect 1650 14500 1850 14600
rect 2350 21200 2550 21300
rect 5750 21300 7350 21500
rect 2350 18200 2400 21200
rect 2500 18200 2550 21200
rect 2350 18000 2550 18200
rect 2650 21200 2950 21250
rect 2650 18200 2700 21200
rect 2900 18200 2950 21200
rect 2650 18150 2950 18200
rect 3050 21200 3250 21250
rect 3050 18200 3100 21200
rect 3200 18200 3250 21200
rect 3050 18000 3250 18200
rect 3750 21200 4550 21250
rect 3750 18200 3800 21200
rect 4500 18200 4550 21200
rect 3750 18150 4550 18200
rect 5050 21200 5250 21250
rect 5050 18200 5100 21200
rect 5200 18200 5250 21200
rect 5050 18000 5250 18200
rect 5350 21200 5650 21250
rect 5350 18200 5400 21200
rect 5600 18200 5650 21200
rect 5350 18150 5650 18200
rect 5750 21200 5950 21300
rect 5750 18200 5800 21200
rect 5900 18200 5950 21200
rect 5750 18000 5950 18200
rect 6450 21200 6650 21250
rect 6450 18200 6500 21200
rect 6600 18200 6650 21200
rect 6450 18100 6650 18200
rect 7150 21200 7350 21300
rect 7150 18200 7200 21200
rect 7300 18200 7350 21200
rect 2350 17800 3250 18000
rect 3300 17950 5000 18000
rect 3300 17850 3350 17950
rect 4950 17850 5000 17950
rect 3300 17800 5000 17850
rect 5050 17800 5950 18000
rect 2350 17600 2550 17800
rect 2350 14600 2400 17600
rect 2500 14600 2550 17600
rect 2350 14550 2550 14600
rect 2650 17600 2950 17650
rect 2650 14600 2700 17600
rect 2900 14600 2950 17600
rect 2650 14550 2950 14600
rect 3050 17600 3250 17800
rect 3050 14600 3100 17600
rect 3200 14600 3250 17600
rect 3050 14550 3250 14600
rect 3750 17600 3950 17650
rect 3750 14600 3800 17600
rect 3900 14600 3950 17600
rect 3750 14550 3950 14600
rect 4350 17600 4550 17650
rect 4350 14600 4400 17600
rect 4500 14600 4550 17600
rect 5050 17600 5250 17800
rect 5050 14600 5100 17600
rect 5200 14600 5250 17600
rect 5350 17600 5650 17650
rect 5350 14600 5400 17600
rect 5600 14600 5650 17600
rect -1150 14450 -100 14500
rect -1150 14350 -450 14450
rect -150 14350 -100 14450
rect -1150 14300 -100 14350
rect 1200 14450 2550 14500
rect 1200 14350 1250 14450
rect 1550 14350 1950 14450
rect 2250 14350 2550 14450
rect 4350 14400 4550 14600
rect 5350 14550 5650 14600
rect 5750 17600 5950 17800
rect 6400 18050 6700 18100
rect 6400 17750 6450 18050
rect 6650 17750 6700 18050
rect 6400 17700 6700 17750
rect 7150 18000 7350 18200
rect 7450 21200 7750 21250
rect 7450 18200 7500 21200
rect 7700 18200 7750 21200
rect 7450 18150 7750 18200
rect 8150 21200 8350 21250
rect 8150 18200 8200 21200
rect 8300 18200 8350 21200
rect 8150 18000 8350 18200
rect 8850 21200 9450 21250
rect 8850 18200 8900 21200
rect 9000 18200 9200 21200
rect 9400 18200 9450 21200
rect 8850 18100 9450 18200
rect 7150 17800 8350 18000
rect 8400 18050 9450 18100
rect 8400 17950 8450 18050
rect 8750 17950 9450 18050
rect 8400 17900 9450 17950
rect 5750 14600 5800 17600
rect 5900 14600 5950 17600
rect 5750 14550 5950 14600
rect 6450 17600 6650 17700
rect 6450 14600 6500 17600
rect 6600 14600 6650 17600
rect 6450 14500 6650 14600
rect 7150 17600 7350 17800
rect 7150 14600 7200 17600
rect 7300 14600 7350 17600
rect 7150 14550 7350 14600
rect 7450 17600 7750 17650
rect 7450 14600 7500 17600
rect 7700 14600 7750 17600
rect 7450 14550 7750 14600
rect 8150 17600 8350 17800
rect 8150 14600 8200 17600
rect 8300 14600 8350 17600
rect 8150 14550 8350 14600
rect 8850 17600 9450 17900
rect 8850 14600 8900 17600
rect 9000 14600 9200 17600
rect 9400 14600 9450 17600
rect 8850 14500 9450 14600
rect 5750 14450 7100 14500
rect 1200 14300 2550 14350
rect 1350 13850 1850 13900
rect 1350 10850 1400 13850
rect 1500 10850 1700 13850
rect 1800 10850 1850 13850
rect 1350 10800 1850 10850
rect 2350 13850 2550 14300
rect 3300 14350 5000 14400
rect 3300 14250 3350 14350
rect 4950 14250 5000 14350
rect 3300 14200 5000 14250
rect 5750 14350 6050 14450
rect 6350 14350 6750 14450
rect 7050 14350 7100 14450
rect 5750 14300 7100 14350
rect 8400 14450 9450 14500
rect 8400 14350 8450 14450
rect 8750 14350 9450 14450
rect 8400 14300 9450 14350
rect 2350 10850 2400 13850
rect 2500 10850 2550 13850
rect 2350 10800 2550 10850
rect 3050 13850 3250 13900
rect 3050 10850 3100 13850
rect 3200 10850 3250 13850
rect 3050 10800 3250 10850
rect 3750 13850 4550 13900
rect 5750 13850 5950 14300
rect 3750 10850 3800 13850
rect 3900 10850 4100 13850
rect 4200 10850 4400 13850
rect 4500 10850 4550 13850
rect 3750 10800 4550 10850
rect 5050 13800 5250 13850
rect 5050 10850 5100 13800
rect 5200 10850 5250 13800
rect 5050 10800 5250 10850
rect 5750 10850 5800 13850
rect 5900 10850 5950 13850
rect 5750 10800 5950 10850
rect 6450 13850 6950 13900
rect 6450 10850 6500 13850
rect 6600 10850 6800 13850
rect 6900 10850 6950 13850
rect 6450 10800 6950 10850
rect 3000 10600 3700 10650
rect 3000 10500 3050 10600
rect 3650 10500 3700 10600
rect 3000 10450 3700 10500
rect 1350 10250 1850 10300
rect 1350 7250 1400 10250
rect 1500 7250 1700 10250
rect 1800 7250 1850 10250
rect 1350 7200 1850 7250
rect 2350 10250 2550 10300
rect 2350 7250 2400 10250
rect 2500 7250 2550 10250
rect 1900 7100 2300 7150
rect 1900 7000 1950 7100
rect 2250 7000 2300 7100
rect 1900 6950 2300 7000
rect 2350 6800 2550 7250
rect 3050 10250 3250 10300
rect 3050 7250 3100 10250
rect 3200 7250 3250 10250
rect 3050 7200 3250 7250
rect 3750 10250 4550 10300
rect 3750 7250 3800 10250
rect 3900 7250 4100 10250
rect 4200 7250 4400 10250
rect 4500 7250 4550 10250
rect 3750 7200 4550 7250
rect 5050 10250 5250 10300
rect 5050 7250 5100 10250
rect 5200 7250 5250 10250
rect 5050 7200 5250 7250
rect 5750 10250 5950 10300
rect 5750 7250 5800 10250
rect 5900 7250 5950 10250
rect -1150 6750 -100 6800
rect -1150 6650 -450 6750
rect -150 6650 -100 6750
rect -1150 6600 -100 6650
rect 1200 6750 2550 6800
rect 1200 6650 1250 6750
rect 1550 6650 1950 6750
rect 2250 6650 2550 6750
rect 3300 6850 5000 6900
rect 3300 6750 3350 6850
rect 4950 6750 5000 6850
rect 3300 6700 5000 6750
rect 5750 6800 5950 7250
rect 6450 10250 6950 10300
rect 6450 7250 6500 10250
rect 6600 7250 6800 10250
rect 6900 7250 6950 10250
rect 6450 7200 6950 7250
rect 6000 7100 6400 7150
rect 6000 7000 6050 7100
rect 6350 7000 6400 7100
rect 6000 6950 6400 7000
rect 9150 6800 9450 14300
rect 5750 6750 7100 6800
rect 1200 6600 2550 6650
rect -1150 6500 -550 6600
rect -1150 3500 -1100 6500
rect -900 3500 -700 6500
rect -600 3500 -550 6500
rect -1150 3200 -550 3500
rect -50 6500 150 6550
rect -50 3500 0 6500
rect 100 3500 150 6500
rect -50 3300 150 3500
rect 550 6500 850 6550
rect 550 3500 600 6500
rect 800 3500 850 6500
rect 550 3450 850 3500
rect 950 6500 1150 6550
rect 950 3500 1000 6500
rect 1100 3500 1150 6500
rect 950 3300 1150 3500
rect 1650 6500 1850 6600
rect 1650 3500 1700 6500
rect 1800 3500 1850 6500
rect 1650 3400 1850 3500
rect 2350 6500 2550 6550
rect 2350 3500 2400 6500
rect 2500 3500 2550 6500
rect -1150 3150 -100 3200
rect -1150 3050 -450 3150
rect -150 3050 -100 3150
rect -1150 3000 -100 3050
rect -50 3100 1150 3300
rect -1150 2900 -550 3000
rect -1150 -100 -1100 2900
rect -900 -100 -700 2900
rect -600 -100 -550 2900
rect -1150 -150 -550 -100
rect -50 2900 150 3100
rect -50 -100 0 2900
rect 100 -100 150 2900
rect -50 -150 150 -100
rect 550 2900 850 2950
rect 550 -100 600 2900
rect 800 -100 850 2900
rect 550 -150 850 -100
rect 950 2900 1150 3100
rect 1600 3350 1900 3400
rect 1600 3050 1650 3350
rect 1850 3050 1900 3350
rect 1600 3000 1900 3050
rect 2350 3300 2550 3500
rect 2650 6500 2950 6550
rect 3750 6500 3950 6700
rect 5750 6650 6050 6750
rect 6350 6650 6750 6750
rect 7050 6650 7100 6750
rect 5750 6600 7100 6650
rect 8400 6750 9450 6800
rect 8400 6650 8450 6750
rect 8750 6650 9450 6750
rect 8400 6600 9450 6650
rect 2650 3500 2700 6500
rect 2900 3500 2950 6500
rect 2650 3450 2950 3500
rect 3050 3500 3100 6500
rect 3200 3500 3250 6500
rect 3050 3300 3250 3500
rect 3750 3500 3800 6500
rect 3900 3500 3950 6500
rect 3750 3450 3950 3500
rect 4350 6500 4550 6550
rect 4350 3500 4400 6500
rect 4500 3500 4550 6500
rect 4350 3450 4550 3500
rect 5050 6500 5250 6550
rect 5050 3500 5100 6500
rect 5200 3500 5250 6500
rect 5050 3300 5250 3500
rect 5350 6500 5650 6550
rect 5350 3500 5400 6500
rect 5600 3500 5650 6500
rect 5350 3450 5650 3500
rect 5750 6500 5950 6550
rect 5750 3500 5800 6500
rect 5900 3500 5950 6500
rect 5750 3300 5950 3500
rect 2350 3100 3250 3300
rect 3300 3250 5000 3300
rect 3300 3150 3350 3250
rect 4950 3150 5000 3250
rect 3300 3100 5000 3150
rect 5050 3100 5950 3300
rect 950 -100 1000 2900
rect 1100 -100 1150 2900
rect 950 -200 1150 -100
rect 1650 2900 1850 3000
rect 1650 -100 1700 2900
rect 1800 -100 1850 2900
rect 1650 -150 1850 -100
rect 2350 2900 2550 3100
rect 2350 -100 2400 2900
rect 2500 -100 2550 2900
rect 2350 -200 2550 -100
rect 2650 2900 2950 2950
rect 2650 -100 2700 2900
rect 2900 -100 2950 2900
rect 2650 -150 2950 -100
rect 3050 2900 3250 3100
rect 3050 -100 3100 2900
rect 3200 -100 3250 2900
rect 3050 -150 3250 -100
rect 3750 2900 4550 2950
rect 3750 -100 3800 2900
rect 4500 -100 4550 2900
rect 3750 -150 4550 -100
rect 5050 2900 5250 3100
rect 5050 -100 5100 2900
rect 5200 -100 5250 2900
rect 5050 -150 5250 -100
rect 5350 2900 5650 2950
rect 5350 -100 5400 2900
rect 5600 -100 5650 2900
rect 5350 -150 5650 -100
rect 5750 2900 5950 3100
rect 5750 -100 5800 2900
rect 5900 -100 5950 2900
rect 5750 -150 5950 -100
rect 6450 6500 6650 6600
rect 6450 3500 6500 6500
rect 6600 3500 6650 6500
rect 6450 2900 6650 3500
rect 6450 -100 6500 2900
rect 6600 -100 6650 2900
rect 6450 -150 6650 -100
rect 7150 6500 7350 6550
rect 7150 3500 7200 6500
rect 7300 3500 7350 6500
rect 7150 3300 7350 3500
rect 7450 6500 7750 6550
rect 7450 3500 7500 6500
rect 7700 3500 7750 6500
rect 7450 3450 7750 3500
rect 8150 6500 8350 6600
rect 8150 3500 8200 6500
rect 8300 3500 8350 6500
rect 8150 3300 8350 3500
rect 7150 3100 8350 3300
rect 8850 6500 9450 6600
rect 8850 3500 8900 6500
rect 9000 3500 9200 6500
rect 9400 3500 9450 6500
rect 8850 3200 9450 3500
rect 7150 2900 7350 3100
rect 7150 -100 7200 2900
rect 7300 -100 7350 2900
rect 7150 -150 7350 -100
rect 7450 2900 7750 2950
rect 7450 -100 7500 2900
rect 7700 -100 7750 2900
rect 7450 -150 7750 -100
rect 8150 2900 8350 3100
rect 8400 3150 9450 3200
rect 8400 3050 8450 3150
rect 8750 3050 9450 3150
rect 8400 3000 9450 3050
rect 8150 -100 8200 2900
rect 8300 -100 8350 2900
rect 8150 -150 8350 -100
rect 8850 2900 9450 3000
rect 8850 -100 8900 2900
rect 9000 -100 9200 2900
rect 9400 -100 9450 2900
rect 8850 -150 9450 -100
rect 950 -400 2550 -200
rect 5800 -300 5900 -150
rect 7200 -300 7300 -150
rect 5800 -400 7300 -300
<< viali >>
rect -1100 18200 -900 21200
rect 600 18200 800 21200
rect -1100 14600 -900 17600
rect 600 14600 800 17600
rect 1000 14600 1100 17600
rect 2700 18200 2900 21200
rect 3800 18200 4500 21200
rect 5400 18200 5600 21200
rect 3350 17850 4950 17950
rect 2700 14600 2900 17600
rect 3800 14600 3900 17600
rect 4400 14600 4500 17600
rect 5400 14600 5600 17600
rect 6450 17750 6650 18050
rect 7500 18200 7700 21200
rect 9200 18200 9400 21200
rect 7200 14600 7300 17600
rect 7500 14600 7700 17600
rect 9200 14600 9400 17600
rect 1400 10850 1500 13850
rect 3350 14250 4250 14350
rect 2400 12700 2500 13850
rect 3100 10850 3200 12100
rect 4100 10850 4200 13850
rect 5100 10850 5200 12100
rect 5800 12700 5900 13850
rect 6800 10850 6900 13850
rect 3050 10500 3650 10600
rect 1400 7250 1500 10250
rect 2400 7250 2500 8400
rect 1950 7000 2250 7100
rect 3100 9000 3200 10250
rect 4100 7250 4200 10250
rect 5100 9000 5200 10250
rect 5800 7250 5900 8400
rect 6800 7250 6900 10250
rect 6050 7000 6350 7100
rect -1100 3500 -900 6500
rect 600 3500 800 6500
rect 1000 3500 1100 6500
rect -1100 -100 -900 2900
rect 600 -100 800 2900
rect 1650 3050 1850 3350
rect 2700 3500 2900 6500
rect 3800 3500 3900 6500
rect 4400 3500 4500 6500
rect 5400 3500 5600 6500
rect 3350 3150 4950 3250
rect 2700 -100 2900 2900
rect 3800 -100 4500 2900
rect 5400 -100 5600 2900
rect 7200 3500 7300 6500
rect 7500 3500 7700 6500
rect 9200 3500 9400 6500
rect 7500 -100 7700 2900
rect 9200 -100 9400 2900
<< metal1 >>
rect -1250 21250 9550 21450
rect -1150 21200 -850 21250
rect -1150 18200 -1100 21200
rect -900 18200 -850 21200
rect -1150 17600 -850 18200
rect -1150 14600 -1100 17600
rect -900 14600 -850 17600
rect -1150 14550 -850 14600
rect 550 21200 850 21250
rect 550 18200 600 21200
rect 800 18200 850 21200
rect 550 17600 850 18200
rect 2650 21200 2950 21250
rect 2650 18200 2700 21200
rect 2900 18200 2950 21200
rect 550 14600 600 17600
rect 800 14600 850 17600
rect 550 14550 850 14600
rect 950 17600 1150 17650
rect 950 14600 1000 17600
rect 1100 14600 1150 17600
rect 950 14550 1150 14600
rect 2650 17600 2950 18200
rect 3750 21200 4550 21250
rect 3750 18200 3800 21200
rect 4500 18200 4550 21200
rect 3750 18150 4550 18200
rect 5350 21200 5650 21250
rect 5350 18200 5400 21200
rect 5600 18200 5650 21200
rect 3300 17950 5000 18000
rect 3300 17850 3350 17950
rect 4950 17850 5000 17950
rect 3300 17800 5000 17850
rect 2650 14600 2700 17600
rect 2900 14600 2950 17600
rect 2650 14550 2950 14600
rect 3750 17600 3950 17650
rect 3750 14600 3800 17600
rect 3900 14600 3950 17600
rect 3750 14550 3950 14600
rect 4350 17600 4550 17650
rect 4350 14600 4400 17600
rect 4500 14600 4550 17600
rect 4350 14550 4550 14600
rect 5350 17600 5650 18200
rect 7450 21200 7750 21250
rect 7450 18200 7500 21200
rect 7700 18200 7750 21200
rect 6400 18050 6700 18100
rect 6400 17750 6450 18050
rect 6650 17750 6700 18050
rect 6400 17700 6700 17750
rect 5350 14600 5400 17600
rect 5600 14600 5650 17600
rect 5350 14550 5650 14600
rect 5750 14550 5950 17650
rect 7150 17600 7350 17650
rect 7150 14600 7200 17600
rect 7300 14600 7350 17600
rect 7150 14550 7350 14600
rect 7450 17600 7750 18200
rect 7450 14600 7500 17600
rect 7700 14600 7750 17600
rect 7450 14550 7750 14600
rect 9150 21200 9450 21250
rect 9150 18200 9200 21200
rect 9400 18200 9450 21200
rect 9150 17600 9450 18200
rect 9150 14600 9200 17600
rect 9400 14600 9450 17600
rect 9150 14550 9450 14600
rect 3300 14350 4300 14400
rect 3300 14250 3350 14350
rect 4250 14250 4300 14350
rect 3300 14200 4300 14250
rect 1350 13850 1550 13900
rect 1350 10850 1400 13850
rect 1500 10850 1550 13850
rect 2350 13850 2550 13900
rect 2350 12700 2400 13850
rect 2500 12700 2550 13850
rect 2350 12650 2550 12700
rect 3750 13850 4550 13900
rect 1350 10250 1550 10850
rect 3050 12100 3250 12150
rect 3050 10850 3100 12100
rect 3200 10850 3250 12100
rect 3050 10800 3250 10850
rect 3750 10850 4100 13850
rect 4200 10850 4550 13850
rect 5750 13850 5950 13900
rect 5750 12700 5800 13850
rect 5900 12700 5950 13850
rect 5750 12650 5950 12700
rect 6750 13850 6950 13900
rect 3750 10800 4550 10850
rect 5050 12100 5250 12150
rect 5050 10850 5100 12100
rect 5200 10850 5250 12100
rect 5050 10800 5250 10850
rect 6750 10850 6800 13850
rect 6900 10850 6950 13850
rect 3000 10600 3700 10650
rect 3000 10500 3050 10600
rect 3650 10500 3700 10600
rect 3000 10450 3700 10500
rect 4050 10300 4250 10800
rect 1350 7250 1400 10250
rect 1500 7250 1550 10250
rect 3050 10250 3250 10300
rect 3050 9000 3100 10250
rect 3200 9000 3250 10250
rect 3050 8950 3250 9000
rect 3750 10250 4550 10300
rect 1350 7150 1550 7250
rect 2350 8400 2550 8450
rect 2350 7250 2400 8400
rect 2500 7250 2550 8400
rect 2350 7200 2550 7250
rect 3750 7250 4100 10250
rect 4200 7250 4550 10250
rect 5050 10250 5250 10300
rect 5050 9000 5100 10250
rect 5200 9000 5250 10250
rect 5050 8950 5250 9000
rect 6750 10250 6950 10850
rect 3750 7200 4550 7250
rect 5750 8400 5950 8450
rect 5750 7250 5800 8400
rect 5900 7250 5950 8400
rect 5750 7200 5950 7250
rect 6750 7250 6800 10250
rect 6900 7250 6950 10250
rect 4050 7150 4250 7200
rect 6750 7150 6950 7250
rect -1250 7100 9550 7150
rect -1250 7000 1950 7100
rect 2250 7000 6050 7100
rect 6350 7000 9550 7100
rect -1250 6950 9550 7000
rect -1150 6500 -850 6550
rect -1150 3500 -1100 6500
rect -900 3500 -850 6500
rect -1150 2900 -850 3500
rect -1150 -100 -1100 2900
rect -900 -100 -850 2900
rect -1150 -150 -850 -100
rect 550 6500 850 6550
rect 550 3500 600 6500
rect 800 3500 850 6500
rect 550 2900 850 3500
rect 950 6500 1150 6550
rect 950 3500 1000 6500
rect 1100 3500 1150 6500
rect 950 3450 1150 3500
rect 2350 3450 2550 6550
rect 2650 6500 2950 6550
rect 2650 3500 2700 6500
rect 2900 3500 2950 6500
rect 1600 3350 1900 3400
rect 1600 3050 1650 3350
rect 1850 3050 1900 3350
rect 1600 3000 1900 3050
rect 550 -100 600 2900
rect 800 -100 850 2900
rect 550 -150 850 -100
rect 2650 2900 2950 3500
rect 3750 6500 3950 6550
rect 3750 3500 3800 6500
rect 3900 3500 3950 6500
rect 3750 3450 3950 3500
rect 4350 6500 4550 6550
rect 4350 3500 4400 6500
rect 4500 3500 4550 6500
rect 4350 3450 4550 3500
rect 5350 6500 5650 6550
rect 5350 3500 5400 6500
rect 5600 3500 5650 6500
rect 3300 3250 5000 3300
rect 3300 3150 3350 3250
rect 4950 3150 5000 3250
rect 3300 3100 5000 3150
rect 2650 -100 2700 2900
rect 2900 -100 2950 2900
rect 2650 -150 2950 -100
rect 3750 2900 4550 2950
rect 3750 -100 3800 2900
rect 4500 -100 4550 2900
rect 3750 -150 4550 -100
rect 5350 2900 5650 3500
rect 7150 6500 7350 6550
rect 7150 3500 7200 6500
rect 7300 3500 7350 6500
rect 7150 3450 7350 3500
rect 7450 6500 7750 6550
rect 7450 3500 7500 6500
rect 7700 3500 7750 6500
rect 5350 -100 5400 2900
rect 5600 -100 5650 2900
rect 5350 -150 5650 -100
rect 7450 2900 7750 3500
rect 7450 -100 7500 2900
rect 7700 -100 7750 2900
rect 7450 -150 7750 -100
rect 9150 6500 9450 6550
rect 9150 3500 9200 6500
rect 9400 3500 9450 6500
rect 9150 2900 9450 3500
rect 9150 -100 9200 2900
rect 9400 -100 9450 2900
rect 9150 -150 9450 -100
rect -1250 -350 9550 -150
<< via1 >>
rect 1000 14600 1100 17600
rect 3350 17850 4950 17950
rect 3800 14600 3900 17600
rect 6450 17750 6650 18050
rect 7200 14600 7300 17600
rect 3350 14250 4250 14350
rect 2400 12700 2500 13850
rect 3100 10850 3200 12100
rect 5800 12700 5900 13850
rect 5100 10850 5200 12100
rect 3050 10500 3650 10600
rect 3100 9000 3200 10250
rect 2400 7250 2500 8400
rect 5100 9000 5200 10250
rect 5800 7250 5900 8400
rect 1000 3500 1100 6500
rect 1650 3050 1850 3350
rect 3800 3500 3900 6500
rect 4400 3500 4500 6500
rect 3350 3150 4950 3250
rect 7200 3500 7300 6500
<< metal2 >>
rect 6400 18050 6700 18100
rect 6400 18000 6450 18050
rect 3300 17950 6450 18000
rect 3300 17850 3350 17950
rect 4950 17850 6450 17950
rect 3300 17800 6450 17850
rect 6400 17750 6450 17800
rect 6650 17750 6700 18050
rect 6400 17700 6700 17750
rect 950 17600 1150 17650
rect 950 14600 1000 17600
rect 1100 14600 1150 17600
rect 950 14550 1150 14600
rect 3750 17600 3950 17650
rect 3750 14600 3800 17600
rect 3900 14750 3950 17600
rect 7150 17600 7350 17650
rect 3900 14600 4550 14750
rect 3750 14550 4550 14600
rect 7150 14600 7200 17600
rect 7300 14600 7350 17600
rect 7150 14550 7350 14600
rect 3300 14350 4300 14400
rect 3300 14250 3350 14350
rect 4250 14250 4300 14350
rect 3300 14200 4300 14250
rect 2350 13850 2550 13900
rect 2350 12700 2400 13850
rect 2500 12700 2550 13850
rect 2350 12650 2550 12700
rect 3750 12600 3950 14200
rect -1250 12200 3950 12600
rect 3050 12100 3250 12150
rect 3050 10850 3100 12100
rect 3200 10850 3250 12100
rect -1250 10650 -850 10850
rect 3050 10800 3250 10850
rect -1250 10600 3700 10650
rect -1250 10500 3050 10600
rect 3650 10500 3700 10600
rect -1250 10450 3700 10500
rect 3050 10250 3250 10300
rect 3050 9000 3100 10250
rect 3200 9000 3250 10250
rect 3050 8950 3250 9000
rect 2350 8400 2550 8450
rect 2350 7250 2400 8400
rect 2500 7250 2550 8400
rect 2350 7200 2550 7250
rect 950 6500 1150 6550
rect 950 3500 1000 6500
rect 1100 3500 1150 6500
rect 950 3450 1150 3500
rect 3750 6500 3950 12200
rect 3750 3500 3800 6500
rect 3900 3500 3950 6500
rect 3750 3450 3950 3500
rect 4350 12600 4550 14550
rect 5750 13850 5950 13900
rect 5750 12700 5800 13850
rect 5900 12700 5950 13850
rect 5750 12650 5950 12700
rect 4350 12200 9550 12600
rect 4350 8900 4550 12200
rect 5050 12100 5250 12150
rect 5050 10850 5100 12100
rect 5200 10850 5250 12100
rect 5050 10800 5250 10850
rect 5050 10250 5250 10300
rect 5050 9000 5100 10250
rect 5200 9000 5250 10250
rect 5050 8950 5250 9000
rect 4350 8500 9550 8900
rect 4350 6500 4550 8500
rect 5750 8400 5950 8450
rect 5750 7250 5800 8400
rect 5900 7250 5950 8400
rect 5750 7200 5950 7250
rect 4350 3500 4400 6500
rect 4500 3500 4550 6500
rect 4350 3450 4550 3500
rect 7150 6500 7350 6550
rect 7150 3500 7200 6500
rect 7300 3500 7350 6500
rect 7150 3450 7350 3500
rect 1600 3350 1900 3400
rect 1600 3050 1650 3350
rect 1850 3300 1900 3350
rect 1850 3250 5000 3300
rect 1850 3150 3350 3250
rect 4950 3150 5000 3250
rect 1850 3100 5000 3150
rect 1850 3050 1900 3100
rect 1600 3000 1900 3050
<< via2 >>
rect 1000 14600 1100 17600
rect 7200 14600 7300 17600
rect 2400 12700 2500 13850
rect 3100 10850 3200 12100
rect 3100 9000 3200 10250
rect 2400 7250 2500 8400
rect 1000 3500 1100 6500
rect 5800 12700 5900 13850
rect 5100 10850 5200 12100
rect 5100 9000 5200 10250
rect 5800 7250 5900 8400
rect 7200 3500 7300 6500
<< metal3 >>
rect 950 17600 1150 17650
rect 950 14750 1000 17600
rect 650 14600 1000 14750
rect 1100 14600 1150 17600
rect 650 14550 1150 14600
rect 7150 17600 7350 17650
rect 7150 14600 7200 17600
rect 7300 14600 7350 17600
rect 650 3350 850 14550
rect 2350 13850 2550 13900
rect 2350 12850 2400 13850
rect 2100 12700 2400 12850
rect 2500 12700 2550 13850
rect 5750 13850 5950 13900
rect 5750 12850 5800 13850
rect 2100 12650 2550 12700
rect 5500 12700 5800 12850
rect 5900 12700 5950 13850
rect 5500 12650 5950 12700
rect 2100 7150 2300 12650
rect 3050 12100 3250 12150
rect 3050 11000 3100 12100
rect 2800 10850 3100 11000
rect 3200 10850 3250 12100
rect 5050 12100 5250 12150
rect 5050 11000 5100 12100
rect 2800 10800 3250 10850
rect 4050 10850 5100 11000
rect 5200 10850 5250 12100
rect 4050 10800 5250 10850
rect 2800 8900 3000 10800
rect 4050 10300 4250 10800
rect 3050 10250 4250 10300
rect 3050 9000 3100 10250
rect 3200 10100 4250 10250
rect 5050 10250 5250 10300
rect 3200 9000 3250 10100
rect 3050 8950 3250 9000
rect 5050 9000 5100 10250
rect 5200 9000 5250 10250
rect 5050 8900 5250 9000
rect 2800 8700 5250 8900
rect 5500 8450 5700 12650
rect 2350 8400 5700 8450
rect 2350 7250 2400 8400
rect 2500 8250 5700 8400
rect 5750 8400 5950 8450
rect 2500 7250 2550 8250
rect 2350 7200 2550 7250
rect 5750 7250 5800 8400
rect 5900 7250 5950 8400
rect 5750 7150 5950 7250
rect 2100 6950 5950 7150
rect 6000 6950 6400 7150
rect 7150 6850 7350 14600
rect 950 6650 7350 6850
rect 950 6500 1150 6650
rect 950 3500 1000 6500
rect 1100 3500 1150 6500
rect 950 3450 1150 3500
rect 7150 6500 7350 6550
rect 7150 3500 7200 6500
rect 7300 3500 7350 6500
rect 7150 3350 7350 3500
rect 650 3150 7350 3350
<< labels >>
flabel metal2 -1250 12400 -1250 12400 0 FreeSans 800 0 0 0 I_IN
port 0 nsew
flabel metal2 -1250 10650 -1250 10650 0 FreeSans 800 0 0 0 VBP
port 1 nsew
flabel metal2 9550 12400 9550 12400 0 FreeSans 800 0 0 0 I_OUT
port 2 nsew
flabel metal1 -1250 7050 -1250 7050 0 FreeSans 800 0 0 0 VP
port 3 nsew
flabel metal1 -1250 -250 -1250 -250 0 FreeSans 800 0 0 0 VN
port 5 nsew
<< end >>
