magic
tech sky130A
timestamp 1701134641
<< error_s >>
rect 16100 6300 16103 6303
rect 16197 6300 16200 6303
rect 16097 6297 16100 6300
rect 16200 6297 16203 6300
rect 16097 6100 16100 6103
rect 16200 6100 16203 6103
rect 16100 6097 16103 6100
rect 16197 6097 16200 6100
<< nmos >>
rect 2600 21900 3000 25100
rect 18300 22000 18700 25200
rect 2600 18300 3000 21500
rect 18100 18300 18500 21500
rect 19600 18300 20000 21500
rect 2600 14500 3000 17700
rect 18100 14500 18500 17700
rect 19600 14500 20000 17700
rect 2600 10900 3000 14100
rect 18300 10800 18700 14000
<< ndiff >>
rect 2300 24900 2600 25100
rect 2300 22100 2400 24900
rect 2500 22100 2600 24900
rect 2300 21900 2600 22100
rect 3000 24900 3300 25100
rect 3000 22100 3100 24900
rect 3200 22100 3300 24900
rect 3000 21900 3300 22100
rect 18000 25000 18300 25200
rect 18000 22200 18100 25000
rect 18200 22200 18300 25000
rect 18000 22000 18300 22200
rect 18700 25000 19000 25200
rect 18700 22200 18800 25000
rect 18900 22200 19000 25000
rect 18700 22000 19000 22200
rect 2300 21300 2600 21500
rect 2300 18500 2400 21300
rect 2500 18500 2600 21300
rect 2300 18300 2600 18500
rect 3000 21300 3300 21500
rect 3000 18500 3100 21300
rect 3200 18500 3300 21300
rect 3000 18300 3300 18500
rect 17800 21300 18100 21500
rect 17800 18500 17900 21300
rect 18000 18500 18100 21300
rect 17800 18300 18100 18500
rect 18500 21300 18800 21500
rect 18500 18500 18600 21300
rect 18700 18500 18800 21300
rect 18500 18300 18800 18500
rect 19300 21300 19600 21500
rect 19300 18500 19400 21300
rect 19500 18500 19600 21300
rect 19300 18300 19600 18500
rect 20000 21300 20300 21500
rect 20000 18500 20100 21300
rect 20200 18500 20300 21300
rect 20000 18300 20300 18500
rect 2300 17500 2600 17700
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 2300 14500 2600 14700
rect 3000 17500 3300 17700
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14500 3300 14700
rect 17800 17500 18100 17700
rect 17800 14700 17900 17500
rect 18000 14700 18100 17500
rect 17800 14500 18100 14700
rect 18500 17500 18800 17700
rect 18500 14700 18600 17500
rect 18700 14700 18800 17500
rect 18500 14500 18800 14700
rect 19300 17500 19600 17700
rect 19300 14700 19400 17500
rect 19500 14700 19600 17500
rect 19300 14500 19600 14700
rect 20000 17500 20300 17700
rect 20000 14700 20100 17500
rect 20200 14700 20300 17500
rect 20000 14500 20300 14700
rect 2300 13900 2600 14100
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 2300 10900 2600 11100
rect 3000 13900 3300 14100
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 10900 3300 11100
rect 18000 13800 18300 14000
rect 18000 11000 18100 13800
rect 18200 11000 18300 13800
rect 18000 10800 18300 11000
rect 18700 13800 19000 14000
rect 18700 11000 18800 13800
rect 18900 11000 19000 13800
rect 18700 10800 19000 11000
<< ndiffc >>
rect 2400 22100 2500 24900
rect 3100 22100 3200 24900
rect 18100 22200 18200 25000
rect 18800 22200 18900 25000
rect 2400 18500 2500 21300
rect 3100 18500 3200 21300
rect 17900 18500 18000 21300
rect 18600 18500 18700 21300
rect 19400 18500 19500 21300
rect 20100 18500 20200 21300
rect 2400 14700 2500 17500
rect 3100 14700 3200 17500
rect 17900 14700 18000 17500
rect 18600 14700 18700 17500
rect 19400 14700 19500 17500
rect 20100 14700 20200 17500
rect 2400 11100 2500 13900
rect 3100 11100 3200 13900
rect 18100 11000 18200 13800
rect 18800 11000 18900 13800
<< psubdiff >>
rect 2000 24900 2300 25100
rect 2000 22100 2100 24900
rect 2200 22100 2300 24900
rect 2000 21900 2300 22100
rect 17700 25000 18000 25200
rect 17700 22200 17800 25000
rect 17900 22200 18000 25000
rect 17700 22000 18000 22200
rect 2000 21300 2300 21500
rect 2000 18500 2100 21300
rect 2200 18500 2300 21300
rect 2000 18300 2300 18500
rect 17530 21400 17800 21500
rect 17530 18400 17600 21400
rect 17700 18400 17800 21400
rect 17530 18300 17800 18400
rect 19000 21300 19300 21500
rect 19000 18500 19100 21300
rect 19200 18500 19300 21300
rect 19000 18300 19300 18500
rect 2000 17500 2300 17700
rect 2000 14700 2100 17500
rect 2200 14700 2300 17500
rect 2000 14500 2300 14700
rect 17530 17600 17800 17700
rect 17530 14600 17600 17600
rect 17700 14600 17800 17600
rect 17530 14500 17800 14600
rect 19000 17500 19300 17700
rect 19000 14700 19100 17500
rect 19200 14700 19300 17500
rect 19000 14500 19300 14700
rect 2000 13900 2300 14100
rect 2000 11100 2100 13900
rect 2200 11100 2300 13900
rect 2000 10900 2300 11100
rect 17700 13800 18000 14000
rect 17700 11000 17800 13800
rect 17900 11000 18000 13800
rect 17700 10800 18000 11000
<< psubdiffcont >>
rect 2100 22100 2200 24900
rect 17800 22200 17900 25000
rect 2100 18500 2200 21300
rect 17600 18400 17700 21400
rect 19100 18500 19200 21300
rect 2100 14700 2200 17500
rect 17600 14600 17700 17600
rect 19100 14700 19200 17500
rect 2100 11100 2200 13900
rect 17800 11000 17900 13800
<< poly >>
rect 18300 25200 18700 25300
rect 2600 25100 3000 25200
rect 18300 21900 18700 22000
rect 2600 21750 3000 21900
rect 2600 21650 2650 21750
rect 2950 21650 3000 21750
rect 18300 21700 20000 21900
rect 2600 21500 3000 21650
rect 18100 21500 18500 21600
rect 19600 21500 20000 21700
rect 2600 17700 3000 18300
rect 18100 18200 18500 18300
rect 19600 18200 20000 18300
rect 17200 18150 18500 18200
rect 17200 17850 18150 18150
rect 18450 17850 18500 18150
rect 17200 17800 18500 17850
rect 19200 18150 20000 18200
rect 19200 17850 19250 18150
rect 19450 17850 20000 18150
rect 19200 17800 20000 17850
rect 18100 17700 18500 17800
rect 19600 17700 20000 17800
rect 2600 14350 3000 14500
rect 18100 14400 18500 14500
rect 2600 14250 2650 14350
rect 2950 14250 3000 14350
rect 19600 14300 20000 14500
rect 2600 14100 3000 14250
rect 18300 14100 20000 14300
rect 18300 14000 18700 14100
rect 2600 10800 3000 10900
rect 18300 10700 18700 10800
<< polycont >>
rect 2650 21650 2950 21750
rect 18150 17850 18450 18150
rect 19250 17850 19450 18150
rect 2650 14250 2950 14350
<< locali >>
rect 17300 25300 18900 25500
rect 17300 25100 17500 25300
rect 18700 25100 18900 25300
rect 17700 25000 18300 25100
rect 2000 24900 2600 25000
rect 2000 22100 2100 24900
rect 2200 22100 2400 24900
rect 2500 22100 2600 24900
rect 2000 22000 2600 22100
rect 3000 24900 3300 25000
rect 3000 22100 3100 24900
rect 3200 22100 3300 24900
rect 17700 22200 17800 25000
rect 17900 22200 18100 25000
rect 18200 22200 18300 25000
rect 17700 22100 18300 22200
rect 18700 25000 19000 25100
rect 18700 22200 18800 25000
rect 18900 22200 19000 25000
rect 18700 22100 19000 22200
rect 3000 22000 3300 22100
rect 2400 21800 2500 22000
rect 17800 21800 17900 22100
rect 2400 21750 3000 21800
rect 2400 21650 2650 21750
rect 2950 21650 3000 21750
rect 2400 21600 3000 21650
rect 17600 21700 17900 21800
rect 2400 21400 2500 21600
rect 17600 21400 17700 21700
rect 18500 21600 20200 21800
rect 18500 21400 18700 21600
rect 20000 21400 20200 21600
rect 2000 21300 2600 21400
rect 2000 18500 2100 21300
rect 2200 18500 2400 21300
rect 2500 18500 2600 21300
rect 2000 18400 2600 18500
rect 3000 21300 3300 21400
rect 3000 18500 3100 21300
rect 3200 18500 3300 21300
rect 3000 18400 3300 18500
rect 17800 21300 18100 21400
rect 17800 18500 17900 21300
rect 18000 18500 18100 21300
rect 17800 18400 18100 18500
rect 18500 21300 18800 21400
rect 18500 18500 18600 21300
rect 18700 18500 18800 21300
rect 18500 18400 18800 18500
rect 19000 21300 19600 21400
rect 19000 18500 19100 21300
rect 19200 18500 19400 21300
rect 19500 18500 19600 21300
rect 19000 18400 19600 18500
rect 20000 21300 20300 21400
rect 20000 18500 20100 21300
rect 20200 18500 20300 21300
rect 20000 18400 20300 18500
rect 2000 17800 3500 18200
rect 17600 17600 17700 18400
rect 18100 18150 18500 18200
rect 18100 17850 18150 18150
rect 18450 17850 18500 18150
rect 18100 17800 18500 17850
rect 19200 18150 19500 18400
rect 19200 17850 19250 18150
rect 19450 17850 19500 18150
rect 19200 17600 19500 17850
rect 2000 17500 2600 17600
rect 2000 14700 2100 17500
rect 2200 14700 2400 17500
rect 2500 14700 2600 17500
rect 2000 14600 2600 14700
rect 3000 17500 3300 17600
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14600 3300 14700
rect 17800 17500 18100 17600
rect 17800 14700 17900 17500
rect 18000 14700 18100 17500
rect 17800 14600 18100 14700
rect 18500 17500 18800 17600
rect 18500 14700 18600 17500
rect 18700 14700 18800 17500
rect 18500 14600 18800 14700
rect 19000 17500 19600 17600
rect 19000 14700 19100 17500
rect 19200 14700 19400 17500
rect 19500 14700 19600 17500
rect 19000 14600 19600 14700
rect 20000 17500 20300 17600
rect 20000 14700 20100 17500
rect 20200 14700 20300 17500
rect 20000 14600 20300 14700
rect 2400 14400 2500 14600
rect 2400 14350 3000 14400
rect 2400 14250 2650 14350
rect 2950 14250 3000 14350
rect 2400 14200 3000 14250
rect 17600 14300 17700 14600
rect 18500 14400 18700 14600
rect 20000 14400 20200 14600
rect 17600 14200 17900 14300
rect 18500 14200 20200 14400
rect 2400 14000 2500 14200
rect 2000 13900 2600 14000
rect 2000 11100 2100 13900
rect 2200 11100 2400 13900
rect 2500 11100 2600 13900
rect 2000 11000 2600 11100
rect 3000 13900 3300 14000
rect 17800 13900 17900 14200
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 11000 3300 11100
rect 17700 13800 18300 13900
rect 17700 11000 17800 13800
rect 17900 11000 18100 13800
rect 18200 11000 18300 13800
rect 17200 10900 17500 11000
rect 17700 10900 18300 11000
rect 18700 13800 19000 13900
rect 18700 11000 18800 13800
rect 18900 11000 19000 13800
rect 18700 10900 19000 11000
rect 17300 10800 17500 10900
rect 18700 10800 18900 10900
rect 17300 10600 18900 10800
<< viali >>
rect 4650 29350 4950 29450
rect 2400 22100 2500 24900
rect 18100 22200 18200 25000
rect 2400 18500 2500 21300
rect 18600 20800 18700 21000
rect 19400 18500 19500 21300
rect 2400 14700 2500 17500
rect 18600 15000 18700 15200
rect 19400 14700 19500 17500
rect 2400 11100 2500 13900
rect 18100 11000 18200 13800
rect 4650 6550 4950 6650
rect 6650 6550 6950 6650
rect 8650 6550 8950 6650
rect 10650 6550 10950 6650
rect 12650 6550 12950 6650
rect 14650 6550 14950 6650
rect 16650 6550 16950 6650
<< metal1 >>
rect 4600 29450 5000 29500
rect 4600 29350 4650 29450
rect 4950 29350 5000 29450
rect 4600 29300 5000 29350
rect 6600 29450 7000 29500
rect 6600 29350 6650 29450
rect 6950 29350 7000 29450
rect 6600 29300 7000 29350
rect 8600 29450 9000 29500
rect 8600 29350 8650 29450
rect 8950 29350 9000 29450
rect 8600 29300 9000 29350
rect 10600 29450 11000 29500
rect 10600 29350 10650 29450
rect 10950 29350 11000 29450
rect 10600 29300 11000 29350
rect 14600 29450 15000 29500
rect 14600 29350 14650 29450
rect 14950 29350 15000 29450
rect 14600 29300 15000 29350
rect 16600 29450 17000 29500
rect 16600 29350 16650 29450
rect 16950 29350 17000 29450
rect 16600 29300 17000 29350
rect 2300 26000 3500 29200
rect 17500 26000 19000 29200
rect 2300 24900 2600 26000
rect 17000 25350 17150 25450
rect 2300 22100 2400 24900
rect 2500 22100 2600 24900
rect 18000 25000 19000 26000
rect 3300 23850 3500 23900
rect 3300 23550 3350 23850
rect 3450 23550 3500 23850
rect 3300 23500 3500 23550
rect 17500 23850 17700 23900
rect 17500 23550 17550 23850
rect 17650 23550 17700 23850
rect 17500 23500 17700 23550
rect 2300 21300 2600 22100
rect 18000 22200 18100 25000
rect 18200 22200 19000 25000
rect 18000 21900 19000 22200
rect 18000 21500 19600 21900
rect 2300 18500 2400 21300
rect 2500 18500 2600 21300
rect 19300 21300 19600 21500
rect 18500 21000 18800 21100
rect 18500 20800 18600 21000
rect 18700 20800 18800 21000
rect 18500 20700 18800 20800
rect 3300 20050 3500 20100
rect 3300 19750 3350 20050
rect 3450 19750 3500 20050
rect 3300 19700 3500 19750
rect 17500 19700 19000 20100
rect 2300 17500 2600 18500
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 18600 16300 19000 19700
rect 19300 18500 19400 21300
rect 19500 18500 19600 21300
rect 19300 18400 19600 18500
rect 3300 16250 3500 16300
rect 3300 15950 3350 16250
rect 3450 15950 3500 16250
rect 3300 15900 3500 15950
rect 17500 15900 19000 16300
rect 19300 17500 19600 17600
rect 18500 15200 18800 15300
rect 18500 15000 18600 15200
rect 18700 15000 18800 15200
rect 18500 14900 18800 15000
rect 2300 13900 2600 14700
rect 19300 14700 19400 17500
rect 19500 14700 19600 17500
rect 19300 14500 19600 14700
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 18000 14100 19600 14500
rect 18000 13800 19000 14100
rect 3300 12450 3500 12500
rect 3300 12150 3350 12450
rect 3450 12150 3500 12450
rect 3300 12100 3500 12150
rect 17500 12450 17700 12500
rect 17500 12150 17550 12450
rect 17650 12150 17700 12450
rect 17500 12100 17700 12150
rect 2300 10000 2600 11100
rect 18000 11000 18100 13800
rect 18200 11000 19000 13800
rect 16950 10550 17150 10650
rect 18000 10000 19000 11000
rect 2300 6800 3500 10000
rect 17500 6800 19000 10000
rect 4600 6650 5000 6700
rect 4600 6550 4650 6650
rect 4950 6550 5000 6650
rect 4600 6500 5000 6550
rect 6600 6650 7000 6700
rect 6600 6550 6650 6650
rect 6950 6550 7000 6650
rect 6600 6500 7000 6550
rect 8600 6650 9000 6700
rect 8600 6550 8650 6650
rect 8950 6550 9000 6650
rect 8600 6500 9000 6550
rect 10600 6650 11000 6700
rect 10600 6550 10650 6650
rect 10950 6550 11000 6650
rect 10600 6500 11000 6550
rect 12600 6650 13000 6700
rect 12600 6550 12650 6650
rect 12950 6550 13000 6650
rect 12600 6500 13000 6550
rect 14600 6650 15000 6700
rect 14600 6550 14650 6650
rect 14950 6550 15000 6650
rect 14600 6500 15000 6550
rect 16600 6650 17000 6700
rect 16600 6550 16650 6650
rect 16950 6550 17000 6650
rect 16600 6500 17000 6550
<< via1 >>
rect 4650 29350 4950 29450
rect 6650 29350 6950 29450
rect 8650 29350 8950 29450
rect 10650 29350 10950 29450
rect 14650 29350 14950 29450
rect 16650 29350 16950 29450
rect 17150 25350 17350 25450
rect 3350 23550 3450 23850
rect 17550 23550 17650 23850
rect 18600 20800 18700 21000
rect 3350 19750 3450 20050
rect 3350 15950 3450 16250
rect 18600 15000 18700 15200
rect 3350 12150 3450 12450
rect 17550 12150 17650 12450
rect 17150 10550 17350 10650
rect 4650 6550 4950 6650
rect 6650 6550 6950 6650
rect 8650 6550 8950 6650
rect 10650 6550 10950 6650
rect 12650 6550 12950 6650
rect 14650 6550 14950 6650
rect 16650 6550 16950 6650
rect 16100 6100 16200 6300
<< metal2 >>
rect 4600 29450 5000 29500
rect 4600 29350 4650 29450
rect 4950 29350 5000 29450
rect 2000 23850 4200 23900
rect 2000 23550 3350 23850
rect 3450 23550 4200 23850
rect 2000 23500 4200 23550
rect 2000 20050 3500 20100
rect 2000 19750 3350 20050
rect 3450 19750 3500 20050
rect 2000 19700 3500 19750
rect 3000 16300 3400 19700
rect 2000 16250 3500 16300
rect 2000 15950 3350 16250
rect 3450 15950 3500 16250
rect 2000 15900 3500 15950
rect 3800 12500 4200 23500
rect 2000 12450 4200 12500
rect 2000 12150 3350 12450
rect 3450 12150 4200 12450
rect 2000 12100 4200 12150
rect 4600 6650 5000 29350
rect 4600 6550 4650 6650
rect 4950 6550 5000 6650
rect 4600 6500 5000 6550
rect 6600 29450 7000 29500
rect 6600 29350 6650 29450
rect 6950 29350 7000 29450
rect 6600 6650 7000 29350
rect 6600 6550 6650 6650
rect 6950 6550 7000 6650
rect 6600 6500 7000 6550
rect 8600 29450 9000 29500
rect 8600 29350 8650 29450
rect 8950 29350 9000 29450
rect 8600 6650 9000 29350
rect 8600 6550 8650 6650
rect 8950 6550 9000 6650
rect 8600 6500 9000 6550
rect 10600 29450 11000 29500
rect 10600 29350 10650 29450
rect 10950 29350 11000 29450
rect 10600 6650 11000 29350
rect 10600 6550 10650 6650
rect 10950 6550 11000 6650
rect 10600 6500 11000 6550
rect 12600 29450 13000 29500
rect 12600 29350 12650 29450
rect 12950 29350 13000 29450
rect 12600 6650 13000 29350
rect 12600 6550 12650 6650
rect 12950 6550 13000 6650
rect 12600 6500 13000 6550
rect 14600 29450 15000 29500
rect 14600 29350 14650 29450
rect 14950 29350 15000 29450
rect 14600 6650 15000 29350
rect 16600 29450 17000 29500
rect 16600 29350 16650 29450
rect 16950 29350 17000 29450
rect 16600 21950 17000 29350
rect 17100 25450 17400 25500
rect 17100 25350 17150 25450
rect 17350 25350 17400 25450
rect 14600 6550 14650 6650
rect 14950 6550 15000 6650
rect 14600 6500 15000 6550
rect 16600 6650 17000 21900
rect 17100 21100 17400 25350
rect 17500 23850 20900 23900
rect 17500 23550 17550 23850
rect 17650 23550 20900 23850
rect 17500 23500 20900 23550
rect 17100 21000 20900 21100
rect 17100 20800 18600 21000
rect 18700 20800 20900 21000
rect 17100 20700 20900 20800
rect 17650 15300 18050 20700
rect 17100 15200 20900 15300
rect 17100 15000 18600 15200
rect 18700 15000 20900 15200
rect 17100 14900 20900 15000
rect 17100 10650 17400 14900
rect 17500 12450 20900 12500
rect 17500 12150 17550 12450
rect 17650 12150 20900 12450
rect 17500 12100 20900 12150
rect 17100 10550 17150 10650
rect 17350 10550 17400 10650
rect 17100 10500 17400 10550
rect 16600 6550 16650 6650
rect 16950 6550 17000 6650
rect 16600 6500 17000 6550
use DAC_block  DAC_block_0
timestamp 1701133304
transform 1 0 13800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_1
timestamp 1701133304
transform 1 0 11800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_2
timestamp 1701133304
transform 1 0 9800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_3
timestamp 1701133304
transform 1 0 7800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_4
timestamp 1701133304
transform 1 0 5800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_5
timestamp 1701133304
transform 1 0 3800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_6
timestamp 1701133304
transform 1 0 1800 0 -1 25300
box 1700 -10800 3700 7300
use DAC_block  DAC_block_14
timestamp 1701133304
transform 1 0 1800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_15
timestamp 1701133304
transform 1 0 13800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_16
timestamp 1701133304
transform 1 0 3800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_17
timestamp 1701133304
transform 1 0 5800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_18
timestamp 1701133304
transform 1 0 7800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_19
timestamp 1701133304
transform 1 0 9800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_20
timestamp 1701133304
transform 1 0 11800 0 1 10700
box 1700 -10800 3700 7300
<< labels >>
flabel metal2 2000 16100 2000 16100 0 FreeSans 800 0 0 0 H_V
port 0 nsew
flabel metal2 2000 19900 2000 19900 0 FreeSans 800 0 0 0 H_V
port 1 nsew
flabel metal2 2000 23700 2000 23700 0 FreeSans 800 0 0 0 I_OUT
port 2 nsew
flabel metal2 2000 12300 2000 12300 0 FreeSans 800 0 0 0 I_OUT
port 3 nsew
flabel locali 2000 18000 2000 18000 0 FreeSans 800 0 0 0 G_V
port 4 nsew
flabel space 4800 -100 4800 -100 0 FreeSans 800 0 0 0 D_6
port 5 nsew
flabel space 6800 -100 6800 -100 0 FreeSans 800 0 0 0 D_5
port 6 nsew
flabel space 8800 -100 8800 -100 0 FreeSans 800 0 0 0 D_4
port 7 nsew
flabel space 10800 -100 10800 -100 0 FreeSans 800 0 0 0 D_3
port 8 nsew
flabel space 12800 -100 12800 -100 0 FreeSans 800 0 0 0 D_2
port 9 nsew
flabel space 14800 -100 14800 -100 0 FreeSans 800 0 0 0 D_1
port 10 nsew
flabel space 16800 -100 16800 -100 0 FreeSans 800 0 0 0 D_0
port 11 nsew
flabel metal2 20900 15100 20900 15100 0 FreeSans 800 0 0 0 I_DUMP
port 12 nsew
flabel metal2 20900 20900 20900 20900 0 FreeSans 800 0 0 0 I_DUMP
port 13 nsew
flabel metal2 20900 12300 20900 12300 0 FreeSans 800 0 0 0 I_OUT_LD
port 14 nsew
flabel metal2 20900 23700 20900 23700 0 FreeSans 800 0 0 0 I_OUT_LD
port 15 nsew
flabel metal1 2300 8300 2300 8300 0 FreeSans 800 0 0 0 VN
port 16 nsew
<< end >>
