magic
tech sky130A
timestamp 1700942202
<< nwell >>
rect -500 -7000 -100 -400
rect 4700 -7000 4900 -400
<< nmos >>
rect 1200 5400 1600 8600
rect 3000 5400 3400 8600
rect 1200 1200 1600 4400
rect 3000 1200 3400 4400
<< ndiff >>
rect -200 8400 1200 8600
rect -200 5600 0 8400
rect 1000 5600 1200 8400
rect -200 5400 1200 5600
rect 1600 8400 3000 8600
rect 1600 5600 1800 8400
rect 2800 5600 3000 8400
rect 1600 5400 3000 5600
rect 3400 8400 4800 8600
rect 3400 5600 3600 8400
rect 4600 5600 4800 8400
rect 3400 5400 4800 5600
rect -200 4200 1200 4400
rect -200 1400 0 4200
rect 1000 1400 1200 4200
rect -200 1200 1200 1400
rect 1600 4200 3000 4400
rect 1600 1400 1800 4200
rect 2800 1400 3000 4200
rect 1600 1200 3000 1400
rect 3400 4200 4800 4400
rect 3400 1400 3600 4200
rect 4600 1400 4800 4200
rect 3400 1200 4800 1400
<< ndiffc >>
rect 0 5600 1000 8400
rect 1800 5600 2800 8400
rect 3600 5600 4600 8400
rect 0 1400 1000 4200
rect 1800 1400 2800 4200
rect 3600 1400 4600 4200
<< poly >>
rect 1200 9050 1600 9100
rect 1200 8750 1250 9050
rect 1550 8750 1600 9050
rect 1200 8600 1600 8750
rect 3000 9050 3400 9100
rect 3000 8750 3050 9050
rect 3350 8750 3400 9050
rect 3000 8600 3400 8750
rect 1200 5300 1600 5400
rect 3000 5300 3400 5400
rect 1200 4400 1600 4500
rect 3000 4400 3400 4500
rect 1200 200 1600 1200
rect 3000 1100 3400 1200
rect 3000 700 4200 1100
rect 1200 -200 3200 200
rect 2800 -500 3200 -200
rect 3800 -50 4200 700
rect 3800 -350 3850 -50
rect 4150 -350 4200 -50
rect 3800 -400 4200 -350
<< polycont >>
rect 1250 8750 1550 9050
rect 3050 8750 3350 9050
rect 3850 -350 4150 -50
<< locali >>
rect -500 9050 4900 9100
rect -500 8750 1250 9050
rect 1550 8750 3050 9050
rect 3350 8750 4900 9050
rect -500 8700 4900 8750
rect -100 8400 1100 8500
rect -100 7200 0 8400
rect -500 6800 0 7200
rect -100 5600 0 6800
rect 1000 5600 1100 8400
rect -100 5500 1100 5600
rect 1700 8400 2900 8500
rect 1700 5600 1800 8400
rect 2800 5600 2900 8400
rect 1700 5500 2900 5600
rect 3500 8400 4700 8500
rect 3500 5600 3600 8400
rect 4600 7200 4700 8400
rect 4600 6800 4900 7200
rect 4600 5600 4700 6800
rect 3500 5500 4700 5600
rect 300 5100 700 5500
rect 300 4700 2500 5100
rect 2100 4300 2500 4700
rect -100 4200 1100 4300
rect -100 2900 0 4200
rect -500 2850 0 2900
rect -500 2550 -450 2850
rect -150 2550 0 2850
rect -500 2500 0 2550
rect -100 1400 0 2500
rect 1000 1400 1100 4200
rect -100 1300 1100 1400
rect 1700 4200 2900 4300
rect 1700 1400 1800 4200
rect 2800 1400 2900 4200
rect 1700 1300 2900 1400
rect 3500 4200 4700 4300
rect 3500 1400 3600 4200
rect 4600 1400 4700 4200
rect 3500 1300 4700 1400
rect 4300 550 4700 1300
rect 4300 250 4350 550
rect 4650 250 4700 550
rect 4300 200 4700 250
rect 3800 -50 4200 0
rect 3800 -350 3850 -50
rect 4150 -350 4200 -50
rect 3800 -500 4200 -350
rect 3700 -600 4200 -500
<< viali >>
rect -450 2550 -150 2850
rect 4350 250 4650 550
<< metal1 >>
rect -500 2850 4900 2900
rect -500 2550 -450 2850
rect -150 2550 4900 2850
rect -500 2500 4900 2550
rect -500 550 4900 600
rect -500 250 4350 550
rect 4650 250 4900 550
rect -500 200 4900 250
rect -500 -6900 -100 -500
rect 4700 -6900 4900 -500
rect -500 -10700 -100 -7500
rect 4700 -10700 4900 -7500
use inverter  inverter_0
timestamp 1700940083
transform 1 0 2500 0 1 -11600
box -2600 800 2200 11200
<< labels >>
rlabel metal1 -500 400 -500 400 7 I_DUMP
port 1 w
rlabel metal1 -500 2700 -500 2700 3 I_OUT
port 2 e
rlabel space 3000 -10800 3000 -10800 5 D_IN
port 3 s
rlabel locali -500 7000 -500 7000 7 H_V
port 5 w
rlabel locali -500 8900 -500 8900 7 G_V
port 4 w
rlabel metal1 -500 -9100 -500 -9100 7 VN
port 6 w
rlabel metal1 -500 -3900 -500 -3900 7 VP
port 7 w
rlabel locali 4900 7000 4900 7000 3 H_V_OUT
port 10 e
rlabel locali 4900 8900 4900 8900 3 G_V_OUT
port 11 e
rlabel metal1 4900 2700 4900 2700 3 I_OUT_OUT
port 9 e
rlabel metal1 4900 400 4900 400 3 I_DUMP_OUT
port 8 e
<< end >>
