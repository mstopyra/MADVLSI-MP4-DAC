magic
tech sky130A
timestamp 1700951739
<< nmos >>
rect -600 24100 -200 27300
rect 40800 24100 41200 27300
rect -600 20000 -200 23200
rect 40600 19900 41000 23100
rect 44000 20000 44400 23200
rect -600 16000 -200 19200
rect 40600 16100 41000 19300
rect 44000 16000 44400 19200
rect -600 11900 -200 15100
rect 40800 11900 41200 15100
<< ndiff >>
rect -2000 27100 -600 27300
rect -2000 24300 -1800 27100
rect -800 24300 -600 27100
rect -2000 24100 -600 24300
rect -200 27100 1200 27300
rect -200 24300 0 27100
rect 1000 24300 1200 27100
rect -200 24100 1200 24300
rect 39400 27100 40800 27300
rect 39400 24300 39600 27100
rect 40600 24300 40800 27100
rect 39400 24100 40800 24300
rect 41200 27100 42600 27300
rect 41200 24300 41400 27100
rect 42400 24300 42600 27100
rect 41200 24100 42600 24300
rect -2000 23000 -600 23200
rect -2000 20200 -1800 23000
rect -800 20200 -600 23000
rect -2000 20000 -600 20200
rect -200 23000 1200 23200
rect -200 20200 0 23000
rect 1000 20200 1200 23000
rect -200 20000 1200 20200
rect 39200 22900 40600 23100
rect 39200 20100 39400 22900
rect 40400 20100 40600 22900
rect 39200 19900 40600 20100
rect 41000 22900 42400 23100
rect 41000 20100 41200 22900
rect 42200 20100 42400 22900
rect 41000 19900 42400 20100
rect 42600 23000 44000 23200
rect 42600 20200 42800 23000
rect 43800 20200 44000 23000
rect 42600 20000 44000 20200
rect 44400 23000 45800 23200
rect 44400 20200 44600 23000
rect 45600 20200 45800 23000
rect 44400 20000 45800 20200
rect -2000 19000 -600 19200
rect -2000 16200 -1800 19000
rect -800 16200 -600 19000
rect -2000 16000 -600 16200
rect -200 19000 1200 19200
rect -200 16200 0 19000
rect 1000 16200 1200 19000
rect -200 16000 1200 16200
rect 39200 19100 40600 19300
rect 39200 16300 39400 19100
rect 40400 16300 40600 19100
rect 39200 16100 40600 16300
rect 41000 19100 42400 19300
rect 41000 16300 41200 19100
rect 42200 16300 42400 19100
rect 41000 16100 42400 16300
rect 42600 19000 44000 19200
rect 42600 16200 42800 19000
rect 43800 16200 44000 19000
rect 42600 16000 44000 16200
rect 44400 19000 45800 19200
rect 44400 16200 44600 19000
rect 45600 16200 45800 19000
rect 44400 16000 45800 16200
rect -2000 14900 -600 15100
rect -2000 12100 -1800 14900
rect -800 12100 -600 14900
rect -2000 11900 -600 12100
rect -200 14900 1200 15100
rect -200 12100 0 14900
rect 1000 12100 1200 14900
rect -200 11900 1200 12100
rect 39400 14900 40800 15100
rect 39400 12100 39600 14900
rect 40600 12100 40800 14900
rect 39400 11900 40800 12100
rect 41200 14900 42600 15100
rect 41200 12100 41400 14900
rect 42400 12100 42600 14900
rect 41200 11900 42600 12100
<< ndiffc >>
rect -1800 24300 -800 27100
rect 0 24300 1000 27100
rect 39600 24300 40600 27100
rect 41400 24300 42400 27100
rect -1800 20200 -800 23000
rect 0 20200 1000 23000
rect 39400 20100 40400 22900
rect 41200 20100 42200 22900
rect 42800 20200 43800 23000
rect 44600 20200 45600 23000
rect -1800 16200 -800 19000
rect 0 16200 1000 19000
rect 39400 16300 40400 19100
rect 41200 16300 42200 19100
rect 42800 16200 43800 19000
rect 44600 16200 45600 19000
rect -1800 12100 -800 14900
rect 0 12100 1000 14900
rect 39600 12100 40600 14900
rect 41400 12100 42400 14900
<< psubdiff >>
rect -3400 27100 -2000 27300
rect -3400 24300 -3200 27100
rect -2200 24300 -2000 27100
rect -3400 24100 -2000 24300
rect 42600 27100 44000 27300
rect 42600 24300 42800 27100
rect 43800 24300 44000 27100
rect 42600 24100 44000 24300
rect -3400 23000 -2000 23200
rect -3400 20200 -3200 23000
rect -2200 20200 -2000 23000
rect -3400 20000 -2000 20200
rect 45800 23000 47200 23200
rect 45800 20200 46000 23000
rect 47000 20200 47200 23000
rect 45800 20000 47200 20200
rect -3400 19000 -2000 19200
rect -3400 16200 -3200 19000
rect -2200 16200 -2000 19000
rect -3400 16000 -2000 16200
rect 45800 19000 47200 19200
rect 45800 16200 46000 19000
rect 47000 16200 47200 19000
rect 45800 16000 47200 16200
rect -3400 14900 -2000 15100
rect -3400 12100 -3200 14900
rect -2200 12100 -2000 14900
rect -3400 11900 -2000 12100
rect 42600 14900 44000 15100
rect 42600 12100 42800 14900
rect 43800 12100 44000 14900
rect 42600 11900 44000 12100
<< psubdiffcont >>
rect -3200 24300 -2200 27100
rect 42800 24300 43800 27100
rect -3200 20200 -2200 23000
rect 46000 20200 47000 23000
rect -3200 16200 -2200 19000
rect 46000 16200 47000 19000
rect -3200 12100 -2200 14900
rect 42800 12100 43800 14900
<< poly >>
rect 10000 32600 10400 32700
rect 10000 32400 10100 32600
rect 10300 32400 10400 32600
rect 10000 32300 10400 32400
rect 15400 32600 15800 32700
rect 15400 32400 15500 32600
rect 15700 32400 15800 32600
rect 15400 32300 15800 32400
rect 20800 32600 21200 32700
rect 20800 32400 20900 32600
rect 21100 32400 21200 32600
rect 20800 32300 21200 32400
rect 26200 32600 26600 32700
rect 26200 32400 26300 32600
rect 26500 32400 26600 32600
rect 26200 32300 26600 32400
rect 31600 32600 32000 32700
rect 31600 32400 31700 32600
rect 31900 32400 32000 32600
rect 31600 32300 32000 32400
rect 37000 32600 37400 32700
rect 37000 32400 37100 32600
rect 37300 32400 37400 32600
rect 37000 32300 37400 32400
rect 40800 27750 41200 27800
rect 40800 27450 40850 27750
rect 41150 27450 41200 27750
rect -600 27300 -200 27400
rect 40800 27300 41200 27450
rect -600 23800 -200 24100
rect 40800 24000 41200 24100
rect -600 23500 -550 23800
rect -250 23500 -200 23800
rect -600 23200 -200 23500
rect 44000 23850 44400 23900
rect 44000 23550 44050 23850
rect 44350 23550 44400 23850
rect 44000 23200 44400 23550
rect 40600 23100 41000 23200
rect -600 19200 -200 20000
rect 44000 19900 44400 20000
rect 40600 19750 41000 19900
rect 40600 19450 40650 19750
rect 40950 19450 41000 19750
rect 40600 19300 41000 19450
rect 44000 19200 44400 19300
rect 40600 16000 41000 16100
rect -600 15700 -200 16000
rect -600 15400 -550 15700
rect -250 15400 -200 15700
rect -600 15100 -200 15400
rect 44000 15650 44400 16000
rect 44000 15350 44050 15650
rect 44350 15350 44400 15650
rect 44000 15300 44400 15350
rect 40800 15100 41200 15200
rect -600 11800 -200 11900
rect 40800 11750 41200 11900
rect 40800 11450 40850 11750
rect 41150 11450 41200 11750
rect 40800 11400 41200 11450
rect 4600 6800 5000 6900
rect 4600 6600 4700 6800
rect 4900 6600 5000 6800
rect 4600 6500 5000 6600
rect 10000 6800 10400 6900
rect 10000 6600 10100 6800
rect 10300 6600 10400 6800
rect 10000 6500 10400 6600
rect 15400 6800 15800 6900
rect 15400 6600 15500 6800
rect 15700 6600 15800 6800
rect 15400 6500 15800 6600
rect 20800 6800 21200 6900
rect 20800 6600 20900 6800
rect 21100 6600 21200 6800
rect 20800 6500 21200 6600
rect 26200 6800 26600 6900
rect 26200 6600 26300 6800
rect 26500 6600 26600 6800
rect 26200 6500 26600 6600
rect 31600 6800 32000 6900
rect 31600 6600 31700 6800
rect 31900 6600 32000 6800
rect 31600 6500 32000 6600
rect 37000 6800 37400 6900
rect 37000 6600 37100 6800
rect 37300 6600 37400 6800
rect 37000 6500 37400 6600
<< polycont >>
rect 10100 32400 10300 32600
rect 15500 32400 15700 32600
rect 20900 32400 21100 32600
rect 26300 32400 26500 32600
rect 31700 32400 31900 32600
rect 37100 32400 37300 32600
rect 40850 27450 41150 27750
rect -550 23500 -250 23800
rect 44050 23550 44350 23850
rect 40650 19450 40950 19750
rect -550 15400 -250 15700
rect 44050 15350 44350 15650
rect 40850 11450 41150 11750
rect 4700 6600 4900 6800
rect 10100 6600 10300 6800
rect 15500 6600 15700 6800
rect 20900 6600 21100 6800
rect 26300 6600 26500 6800
rect 31700 6600 31900 6800
rect 37100 6600 37300 6800
<< locali >>
rect 10000 32650 10400 32700
rect 10000 32350 10050 32650
rect 10350 32350 10400 32650
rect 10000 32300 10400 32350
rect 15400 32650 15800 32700
rect 15400 32350 15450 32650
rect 15750 32350 15800 32650
rect 15400 32300 15800 32350
rect 20800 32650 21200 32700
rect 20800 32350 20850 32650
rect 21150 32350 21200 32650
rect 20800 32300 21200 32350
rect 26200 32650 26600 32700
rect 26200 32350 26250 32650
rect 26550 32350 26600 32650
rect 26200 32300 26600 32350
rect 31600 32650 32000 32700
rect 31600 32350 31650 32650
rect 31950 32350 32000 32650
rect 31600 32300 32000 32350
rect 37000 32650 37400 32700
rect 37000 32350 37050 32650
rect 37350 32350 37400 32650
rect 37000 32300 37400 32350
rect 40800 27750 41700 27800
rect 40800 27450 40850 27750
rect 41150 27450 41700 27750
rect 40800 27400 41700 27450
rect 41300 27200 41700 27400
rect -3300 27100 -700 27200
rect -3300 24300 -3200 27100
rect -2200 24300 -1800 27100
rect -800 24300 -700 27100
rect -3300 24200 -700 24300
rect -100 27100 1100 27200
rect -100 24300 0 27100
rect 1000 26000 1100 27100
rect 39500 27100 40700 27200
rect 39500 26000 39600 27100
rect 1000 25600 1300 26000
rect 39400 25600 39600 26000
rect 1000 24300 1100 25600
rect 39500 24600 39600 25600
rect -100 24200 1100 24300
rect 38900 24300 39600 24600
rect 40600 24300 40700 27100
rect 38900 24200 40700 24300
rect 41300 27100 43900 27200
rect 41300 24300 41400 27100
rect 42400 24300 42800 27100
rect 43800 24600 43900 27100
rect 43800 24300 44400 24600
rect 41300 24200 44400 24300
rect -1150 23850 -700 24200
rect 44000 23900 44400 24200
rect 44000 23850 44900 23900
rect -1150 23800 -200 23850
rect -1150 23500 -550 23800
rect -250 23500 -200 23800
rect 44000 23550 44050 23850
rect 44350 23550 44900 23850
rect 44000 23500 44900 23550
rect -1150 23450 -200 23500
rect 41900 23450 42300 23500
rect -1150 23100 -700 23450
rect 41900 23150 41950 23450
rect 42250 23150 42300 23450
rect -3300 23000 -700 23100
rect -3300 20200 -3200 23000
rect -2200 20200 -1800 23000
rect -800 20200 -700 23000
rect -3300 20100 -700 20200
rect -100 23000 1100 23100
rect 41900 23000 42300 23150
rect 44500 23100 44900 23500
rect -100 20200 0 23000
rect 1000 21700 1100 23000
rect 39300 22900 40500 23000
rect 39300 21700 39400 22900
rect 1000 21650 1300 21700
rect 1000 21350 1250 21650
rect 1000 21300 1300 21350
rect 39100 21300 39400 21700
rect 1000 20200 1100 21300
rect -100 20100 1100 20200
rect 39300 20100 39400 21300
rect 40400 20100 40500 22900
rect 39300 20000 40500 20100
rect 41100 22900 42300 23000
rect 41100 20100 41200 22900
rect 42200 21700 42300 22900
rect 42700 23000 43900 23100
rect 42700 21700 42800 23000
rect 42200 21300 42800 21700
rect 42200 20100 42300 21300
rect 42700 20200 42800 21300
rect 43800 20200 43900 23000
rect 42700 20100 43900 20200
rect 44500 23000 47100 23100
rect 44500 20200 44600 23000
rect 45600 20200 46000 23000
rect 47000 20200 47100 23000
rect 44500 20100 47100 20200
rect 41100 20000 42300 20100
rect -4100 19400 1300 19800
rect 39100 19750 41000 19800
rect 39100 19450 40650 19750
rect 40950 19450 41000 19750
rect 39100 19400 41000 19450
rect 39300 19100 40500 19200
rect -3300 19000 -700 19100
rect -3300 16200 -3200 19000
rect -2200 16200 -1800 19000
rect -800 16200 -700 19000
rect -3300 16100 -700 16200
rect -100 19000 1100 19100
rect -100 16200 0 19000
rect 1000 17900 1100 19000
rect 39300 17900 39400 19100
rect 1000 17850 1300 17900
rect 1000 17550 1250 17850
rect 1000 17500 1300 17550
rect 39100 17500 39400 17900
rect 1000 16200 1100 17500
rect 39300 16300 39400 17500
rect 40400 16300 40500 19100
rect 39300 16200 40500 16300
rect 41100 19100 42300 19200
rect 41100 16300 41200 19100
rect 42200 17900 42300 19100
rect 42700 19000 43900 19100
rect 42700 17900 42800 19000
rect 42200 17500 42800 17900
rect 42200 16300 42300 17500
rect 41100 16200 42300 16300
rect -100 16100 1100 16200
rect -1150 15750 -700 16100
rect 41900 16050 42300 16200
rect 42700 16200 42800 17500
rect 43800 16200 43900 19000
rect 42700 16100 43900 16200
rect 44500 19000 47100 19100
rect 44500 16200 44600 19000
rect 45600 16200 46000 19000
rect 47000 16200 47100 19000
rect 44500 16100 47100 16200
rect 41900 15750 41950 16050
rect 42250 15750 42300 16050
rect -1150 15700 -200 15750
rect 41900 15700 42300 15750
rect 44500 15700 44900 16100
rect -1150 15400 -550 15700
rect -250 15400 -200 15700
rect -1150 15350 -200 15400
rect 44000 15650 44900 15700
rect 44000 15350 44050 15650
rect 44350 15350 44900 15650
rect -1150 15000 -700 15350
rect 44000 15300 44900 15350
rect 44000 15000 44400 15300
rect -3300 14900 -700 15000
rect -3300 12100 -3200 14900
rect -2200 12100 -1800 14900
rect -800 12100 -700 14900
rect -3300 12000 -700 12100
rect -100 14900 1100 15000
rect -100 12100 0 14900
rect 1000 13600 1100 14900
rect 38900 14900 40700 15000
rect 38900 14600 39600 14900
rect 39500 13600 39600 14600
rect 1000 13200 1300 13600
rect 39400 13200 39600 13600
rect 1000 12100 1100 13200
rect -100 12000 1100 12100
rect 39500 12100 39600 13200
rect 40600 12100 40700 14900
rect 39500 12000 40700 12100
rect 41300 14900 44400 15000
rect 41300 12100 41400 14900
rect 42400 12100 42800 14900
rect 43800 14600 44400 14900
rect 43800 12100 43900 14600
rect 41300 12000 43900 12100
rect 41300 11800 41700 12000
rect 40800 11750 41700 11800
rect 40800 11450 40850 11750
rect 41150 11450 41700 11750
rect 40800 11400 41700 11450
rect 4600 6850 5000 6900
rect 4600 6550 4650 6850
rect 4950 6550 5000 6850
rect 4600 6500 5000 6550
rect 10000 6850 10400 6900
rect 10000 6550 10050 6850
rect 10350 6550 10400 6850
rect 10000 6500 10400 6550
rect 15400 6850 15800 6900
rect 15400 6550 15450 6850
rect 15750 6550 15800 6850
rect 15400 6500 15800 6550
rect 20800 6850 21200 6900
rect 20800 6550 20850 6850
rect 21150 6550 21200 6850
rect 20800 6500 21200 6550
rect 26200 6850 26600 6900
rect 26200 6550 26250 6850
rect 26550 6550 26600 6850
rect 26200 6500 26600 6550
rect 31600 6850 32000 6900
rect 31600 6550 31650 6850
rect 31950 6550 32000 6850
rect 31600 6500 32000 6550
rect 37000 6850 37400 6900
rect 37000 6550 37050 6850
rect 37350 6550 37400 6850
rect 37000 6500 37400 6550
<< viali >>
rect 4650 32350 4950 32650
rect 10050 32600 10350 32650
rect 10050 32400 10100 32600
rect 10100 32400 10300 32600
rect 10300 32400 10350 32600
rect 10050 32350 10350 32400
rect 15450 32600 15750 32650
rect 15450 32400 15500 32600
rect 15500 32400 15700 32600
rect 15700 32400 15750 32600
rect 15450 32350 15750 32400
rect 20850 32600 21150 32650
rect 20850 32400 20900 32600
rect 20900 32400 21100 32600
rect 21100 32400 21150 32600
rect 20850 32350 21150 32400
rect 26250 32600 26550 32650
rect 26250 32400 26300 32600
rect 26300 32400 26500 32600
rect 26500 32400 26550 32600
rect 26250 32350 26550 32400
rect 31650 32600 31950 32650
rect 31650 32400 31700 32600
rect 31700 32400 31900 32600
rect 31900 32400 31950 32600
rect 31650 32350 31950 32400
rect 37050 32600 37350 32650
rect 37050 32400 37100 32600
rect 37100 32400 37300 32600
rect 37300 32400 37350 32600
rect 37050 32350 37350 32400
rect 1350 27950 1650 28250
rect -1800 24300 -800 27100
rect 41400 24300 42400 27100
rect 41950 23150 42250 23450
rect -1800 20200 -800 23000
rect 1250 21350 1550 21650
rect 44600 20200 45600 23000
rect -1800 16200 -800 19000
rect 1250 17550 1550 17850
rect 44600 16200 45600 19000
rect 41950 15750 42250 16050
rect -1800 12100 -800 14900
rect 41400 12100 42400 14900
rect 4650 6800 4950 6850
rect 4650 6600 4700 6800
rect 4700 6600 4900 6800
rect 4900 6600 4950 6800
rect 4650 6550 4950 6600
rect 10050 6800 10350 6850
rect 10050 6600 10100 6800
rect 10100 6600 10300 6800
rect 10300 6600 10350 6800
rect 10050 6550 10350 6600
rect 15450 6800 15750 6850
rect 15450 6600 15500 6800
rect 15500 6600 15700 6800
rect 15700 6600 15750 6800
rect 15450 6550 15750 6600
rect 20850 6800 21150 6850
rect 20850 6600 20900 6800
rect 20900 6600 21100 6800
rect 21100 6600 21150 6800
rect 20850 6550 21150 6600
rect 26250 6800 26550 6850
rect 26250 6600 26300 6800
rect 26300 6600 26500 6800
rect 26500 6600 26550 6800
rect 26250 6550 26550 6600
rect 31650 6800 31950 6850
rect 31650 6600 31700 6800
rect 31700 6600 31900 6800
rect 31900 6600 31950 6800
rect 31650 6550 31950 6600
rect 37050 6800 37350 6850
rect 37050 6600 37100 6800
rect 37100 6600 37300 6800
rect 37300 6600 37350 6800
rect 37050 6550 37350 6600
<< metal1 >>
rect 4600 32650 5000 32700
rect 4600 32350 4650 32650
rect 4950 32350 5000 32650
rect 4600 32300 5000 32350
rect 10000 32650 10400 32700
rect 10000 32350 10050 32650
rect 10350 32350 10400 32650
rect 10000 32300 10400 32350
rect 15400 32650 15800 32700
rect 15400 32350 15450 32650
rect 15750 32350 15800 32650
rect 15400 32300 15800 32350
rect 20800 32650 21200 32700
rect 20800 32350 20850 32650
rect 21150 32350 21200 32650
rect 20800 32300 21200 32350
rect 26200 32650 26600 32700
rect 26200 32350 26250 32650
rect 26550 32350 26600 32650
rect 26200 32300 26600 32350
rect 31600 32650 32000 32700
rect 31600 32350 31650 32650
rect 31950 32350 32000 32650
rect 31600 32300 32000 32350
rect 37000 32650 37400 32700
rect 37000 32350 37050 32650
rect 37350 32350 37400 32650
rect 37000 32300 37400 32350
rect -2000 29000 2000 32200
rect 39100 29000 42600 32200
rect -2000 27100 -600 29000
rect -2000 24300 -1800 27100
rect -800 24300 -600 27100
rect 41200 27100 42600 29000
rect 39000 25950 39400 26000
rect 39000 25650 39050 25950
rect 39350 25650 39400 25950
rect 39000 25600 39400 25650
rect -2000 23000 -600 24300
rect 41200 24300 41400 27100
rect 42400 24300 42600 27100
rect 41200 24100 42600 24300
rect 41900 23450 42300 23500
rect 41900 23150 41950 23450
rect 42250 23150 42300 23450
rect 41900 23100 42300 23150
rect -2000 20200 -1800 23000
rect -800 20200 -600 23000
rect 44400 23000 45800 23200
rect 1200 21650 1600 21700
rect 1200 21350 1250 21650
rect 1550 21350 1600 21650
rect 1200 21300 1600 21350
rect -2000 19000 -600 20200
rect -2000 16200 -1800 19000
rect -800 16200 -600 19000
rect 44400 20200 44600 23000
rect 45600 20200 45800 23000
rect 44400 19000 45800 20200
rect 1200 17850 1600 17900
rect 1200 17550 1250 17850
rect 1550 17550 1600 17850
rect 1200 17500 1600 17550
rect -2000 14900 -600 16200
rect 44400 16200 44600 19000
rect 45600 16200 45800 19000
rect 41900 16050 42300 16100
rect 41900 15750 41950 16050
rect 42250 15750 42300 16050
rect 44400 16000 45800 16200
rect 41900 15700 42300 15750
rect -2000 12100 -1800 14900
rect -800 12100 -600 14900
rect 41200 14900 42600 15100
rect 39000 13550 39400 13600
rect 39000 13250 39050 13550
rect 39350 13250 39400 13550
rect 39000 13200 39400 13250
rect -2000 10200 -600 12100
rect 41200 12100 41400 14900
rect 42400 12100 42600 14900
rect 41200 10200 42600 12100
rect -2000 7000 1700 10200
rect 39100 7000 42600 10200
rect 4600 6850 5000 6900
rect 4600 6550 4650 6850
rect 4950 6550 5000 6850
rect 4600 6500 5000 6550
rect 10000 6850 10400 6900
rect 10000 6550 10050 6850
rect 10350 6550 10400 6850
rect 10000 6500 10400 6550
rect 15400 6850 15800 6900
rect 15400 6550 15450 6850
rect 15750 6550 15800 6850
rect 15400 6500 15800 6550
rect 20800 6850 21200 6900
rect 20800 6550 20850 6850
rect 21150 6550 21200 6850
rect 20800 6500 21200 6550
rect 26200 6850 26600 6900
rect 26200 6550 26250 6850
rect 26550 6550 26600 6850
rect 26200 6500 26600 6550
rect 31600 6850 32000 6900
rect 31600 6550 31650 6850
rect 31950 6550 32000 6850
rect 31600 6500 32000 6550
rect 37000 6850 37400 6900
rect 37000 6550 37050 6850
rect 37350 6550 37400 6850
rect 37000 6500 37400 6550
<< via1 >>
rect 4650 32350 4950 32650
rect 10050 32350 10350 32650
rect 15450 32350 15750 32650
rect 20850 32350 21150 32650
rect 26250 32350 26550 32650
rect 31650 32350 31950 32650
rect 37050 32350 37350 32650
rect 1350 27950 1650 28250
rect 38550 27950 38850 28250
rect 1350 25650 1650 25950
rect 39050 25650 39350 25950
rect 41950 23150 42250 23450
rect 1250 21350 1550 21650
rect 1250 17550 1550 17850
rect 41950 15750 42250 16050
rect 1350 13250 1650 13550
rect 39050 13250 39350 13550
rect 1350 10950 1650 11250
rect 38550 10950 38850 11250
rect 4650 6550 4950 6850
rect 10050 6550 10350 6850
rect 15450 6550 15750 6850
rect 20850 6550 21150 6850
rect 26250 6550 26550 6850
rect 31650 6550 31950 6850
rect 37050 6550 37350 6850
<< metal2 >>
rect 4600 32650 5000 32700
rect 4600 32350 4650 32650
rect 4950 32350 5000 32650
rect -4100 28250 3400 28300
rect -4100 27950 1350 28250
rect 1650 27950 3400 28250
rect -4100 27900 3400 27950
rect -4100 25950 2500 26000
rect -4100 25650 1350 25950
rect 1650 25650 2500 25950
rect -4100 25600 2500 25650
rect -4100 21650 1600 21700
rect -4100 21350 1250 21650
rect 1550 21350 1600 21650
rect -4100 21300 1600 21350
rect 1200 17900 1600 21300
rect -4100 17850 1600 17900
rect -4100 17550 1250 17850
rect 1550 17550 1600 17850
rect -4100 17500 1600 17550
rect 2100 13600 2500 25600
rect -4100 13550 2500 13600
rect -4100 13250 1350 13550
rect 1650 13250 2500 13550
rect -4100 13200 2500 13250
rect 3000 11300 3400 27900
rect -4100 11250 3400 11300
rect -4100 10950 1350 11250
rect 1650 10950 3400 11250
rect -4100 10900 3400 10950
rect 4600 6850 5000 32350
rect 4600 6550 4650 6850
rect 4950 6550 5000 6850
rect 4600 6500 5000 6550
rect 10000 32650 10400 32700
rect 10000 32350 10050 32650
rect 10350 32350 10400 32650
rect 10000 6850 10400 32350
rect 10000 6550 10050 6850
rect 10350 6550 10400 6850
rect 10000 6500 10400 6550
rect 15400 32650 15800 32700
rect 15400 32350 15450 32650
rect 15750 32350 15800 32650
rect 15400 6850 15800 32350
rect 15400 6550 15450 6850
rect 15750 6550 15800 6850
rect 15400 6500 15800 6550
rect 20800 32650 21200 32700
rect 20800 32350 20850 32650
rect 21150 32350 21200 32650
rect 20800 6850 21200 32350
rect 20800 6550 20850 6850
rect 21150 6550 21200 6850
rect 20800 6500 21200 6550
rect 26200 32650 26600 32700
rect 26200 32350 26250 32650
rect 26550 32350 26600 32650
rect 26200 6850 26600 32350
rect 26200 6550 26250 6850
rect 26550 6550 26600 6850
rect 26200 6500 26600 6550
rect 31600 32650 32000 32700
rect 31600 32350 31650 32650
rect 31950 32350 32000 32650
rect 31600 6850 32000 32350
rect 31600 6550 31650 6850
rect 31950 6550 32000 6850
rect 31600 6500 32000 6550
rect 37000 32650 37400 32700
rect 37000 32350 37050 32650
rect 37350 32350 37400 32650
rect 37000 6850 37400 32350
rect 38100 28250 44700 28300
rect 38100 27950 38550 28250
rect 38850 27950 44700 28250
rect 38100 27900 44700 27950
rect 38100 23800 38500 27900
rect 39000 25950 44700 26000
rect 39000 25650 39050 25950
rect 39350 25650 44700 25950
rect 39000 25600 44700 25650
rect 38100 23450 42300 23800
rect 38100 23400 41950 23450
rect 38100 15800 38500 23400
rect 41900 23150 41950 23400
rect 42250 23150 42300 23450
rect 41900 23100 42300 23150
rect 41900 16050 42300 16100
rect 41900 15800 41950 16050
rect 38100 15750 41950 15800
rect 42250 15750 42300 16050
rect 38100 15400 42300 15750
rect 38100 11300 38500 15400
rect 43400 13600 43800 25600
rect 39000 13550 44700 13600
rect 39000 13250 39050 13550
rect 39350 13250 44700 13550
rect 39000 13200 44700 13250
rect 38100 11250 44700 11300
rect 38100 10950 38550 11250
rect 38850 10950 44700 11250
rect 38100 10900 44700 10950
rect 37000 6550 37050 6850
rect 37350 6550 37400 6850
rect 37000 6500 37400 6550
use DAC_block  DAC_block_0
timestamp 1700946606
transform 1 0 34200 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_1
timestamp 1700946606
transform 1 0 1800 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_2
timestamp 1700946606
transform 1 0 7200 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_3
timestamp 1700946606
transform 1 0 12600 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_4
timestamp 1700946606
transform 1 0 18000 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_5
timestamp 1700946606
transform 1 0 23400 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_6
timestamp 1700946606
transform 1 0 28800 0 -1 28500
box -500 -10800 4900 9100
use DAC_block  DAC_block_7
timestamp 1700946606
transform 1 0 34200 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_8
timestamp 1700946606
transform 1 0 28800 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_9
timestamp 1700946606
transform 1 0 23400 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_10
timestamp 1700946606
transform 1 0 18000 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_11
timestamp 1700946606
transform 1 0 12600 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_12
timestamp 1700946606
transform 1 0 7200 0 1 10700
box -500 -10800 4900 9100
use DAC_block  DAC_block_13
timestamp 1700946606
transform 1 0 1800 0 1 10700
box -500 -10800 4900 9100
<< labels >>
rlabel locali 1300 13400 1300 13400 7 H_V
port 5 w
rlabel viali 1300 17700 1300 17700 3 I_OUT
port 2 e
<< end >>
