magic
tech sky130A
timestamp 1701144897
<< error_p >>
rect 3400 3800 3700 7000
rect 3400 1366 3700 3300
<< nwell >>
rect 1700 -10800 2100 -4200
rect 3500 -10800 3700 -4200
<< nmos >>
rect 2300 3800 2700 7000
rect 3000 3800 3400 7000
rect 2300 100 2700 3300
rect 3000 100 3400 3300
<< ndiff >>
rect 2000 6800 2300 7000
rect 2000 4000 2100 6800
rect 2200 4000 2300 6800
rect 2000 3800 2300 4000
rect 2700 6800 3000 7000
rect 2700 4000 2800 6800
rect 2900 4000 3000 6800
rect 2700 3800 3000 4000
rect 3400 6800 3700 7000
rect 3400 4000 3500 6800
rect 3600 4000 3700 6800
rect 3400 3800 3700 4000
rect 2000 3100 2300 3300
rect 2000 300 2100 3100
rect 2200 300 2300 3100
rect 2000 100 2300 300
rect 2700 3100 3000 3300
rect 2700 300 2800 3100
rect 2900 300 3000 3100
rect 2700 100 3000 300
rect 3400 3100 3700 3300
rect 3400 300 3500 3100
rect 3600 300 3700 3100
rect 3400 100 3700 300
<< ndiffc >>
rect 2100 4000 2200 6800
rect 2800 4000 2900 6800
rect 3500 4000 3600 6800
rect 2100 300 2200 3100
rect 2800 300 2900 3100
rect 3500 300 3600 3100
<< psubdiff >>
rect 1700 6900 2000 7000
rect 1700 3900 1800 6900
rect 1900 3900 2000 6900
rect 1700 3800 2000 3900
rect 1700 3200 2000 3300
rect 1700 200 1800 3200
rect 1900 200 2000 3200
rect 1700 100 2000 200
<< psubdiffcont >>
rect 1800 3900 1900 6900
rect 1800 200 1900 3200
<< poly >>
rect 2300 7250 2700 7300
rect 2300 7150 2350 7250
rect 2650 7150 2700 7250
rect 2300 7000 2700 7150
rect 3000 7250 3400 7300
rect 3000 7150 3050 7250
rect 3350 7150 3400 7250
rect 3000 7000 3400 7150
rect 2300 3700 2700 3800
rect 3000 3700 3400 3800
rect 2300 3300 2700 3400
rect 3000 3300 3400 3400
rect 2300 -400 2700 100
rect 3000 -50 3400 100
rect 3000 -150 3050 -50
rect 3350 -150 3400 -50
rect 3000 -200 3400 -150
rect 2300 -600 3200 -400
<< polycont >>
rect 2350 7150 2650 7250
rect 3050 7150 3350 7250
rect 3050 -150 3350 -50
<< locali >>
rect 1700 7250 3700 7300
rect 1700 7150 2350 7250
rect 2650 7150 3050 7250
rect 3350 7150 3700 7250
rect 1700 7100 3700 7150
rect 1800 6900 1900 7000
rect 2000 6800 2300 6900
rect 2000 4000 2100 6800
rect 2200 4000 2300 6800
rect 2000 3900 2300 4000
rect 2700 6800 3000 6900
rect 2700 4000 2800 6800
rect 2900 4000 3000 6800
rect 2700 3900 3000 4000
rect 3400 6800 3700 6900
rect 3400 4000 3500 6800
rect 3600 4000 3700 6800
rect 3400 3900 3700 4000
rect 1800 3200 1900 3900
rect 2100 3600 2200 3900
rect 2100 3500 2900 3600
rect 2800 3200 2900 3500
rect 2000 3100 2300 3200
rect 2000 300 2100 3100
rect 2200 300 2300 3100
rect 2000 200 2300 300
rect 2700 3100 3000 3200
rect 2700 300 2800 3100
rect 2900 300 3000 3100
rect 2700 200 3000 300
rect 3400 3100 3700 3200
rect 3400 300 3500 3100
rect 3600 300 3700 3100
rect 3400 200 3700 300
rect 1800 -700 1900 200
rect 3500 0 3600 200
rect 3000 -50 3400 0
rect 3000 -150 3050 -50
rect 3350 -150 3400 -50
rect 3000 -200 3400 -150
rect 3450 -50 3650 0
rect 3450 -150 3500 -50
rect 3600 -150 3650 -50
rect 3450 -200 3650 -150
rect 3300 -700 3400 -200
rect 1800 -800 2200 -700
<< viali >>
rect 2100 5300 2200 5500
rect 3500 5300 3600 5500
rect 2100 1500 2200 1700
rect 3500 -150 3600 -50
<< metal1 >>
rect 1700 5500 2300 5600
rect 1700 5300 2100 5500
rect 2200 5300 2300 5500
rect 1700 5200 2300 5300
rect 3400 5500 3700 5600
rect 3400 5300 3500 5500
rect 3600 5300 3700 5500
rect 3400 5200 3700 5300
rect 1700 1700 3700 1800
rect 1700 1500 2100 1700
rect 2200 1500 3700 1700
rect 1700 1400 3700 1500
rect 1700 -50 3700 0
rect 1700 -150 3500 -50
rect 3600 -150 3700 -50
rect 1700 -200 3700 -150
rect 1700 -3900 2100 -700
rect 3500 -3900 3700 -700
rect 1700 -10700 2100 -4300
rect 3500 -10700 3700 -4300
use inverter  inverter_0
timestamp 1701117479
transform 1 0 2500 0 1 -11600
box -400 800 1100 11000
<< labels >>
rlabel metal1 1700 -7300 1700 -7300 7 VP
port 7 w
rlabel metal1 1700 -2300 1700 -2300 7 VN
port 6 w
rlabel metal1 1700 1600 1700 1600 3 I_OUT
port 2 e
rlabel metal1 1700 5400 1700 5400 7 H_V
port 5 w
rlabel poly 3000 -600 3000 -600 1 D_IN
port 3 s
rlabel metal1 3700 -50 3700 -50 3 I_DUMP_OUT
port 8 e
rlabel metal1 3700 1650 3700 1650 3 I_OUT_OUT
port 9 e
rlabel locali 3700 7250 3700 7250 3 G_V_OUT
port 11 e
rlabel metal1 3700 5450 3700 5450 3 H_V_OUT
port 10 e
rlabel metal1 1700 -50 1700 -50 7 I_DUMP
port 1 w
<< end >>
