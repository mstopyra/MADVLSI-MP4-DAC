magic
tech sky130A
timestamp 1701123401
<< error_p >>
rect 1500 10897 1600 10900
rect 1500 7903 1503 10897
rect 1597 7903 1600 10897
rect 1500 7900 1600 7903
rect -100 3096 0 3100
<< nmos >>
rect 2000 7800 2400 11000
rect 2700 7800 3100 11000
rect 4900 7800 5300 11000
rect 5600 7800 6000 11000
rect 7500 7800 7900 11000
rect 2800 3900 3200 7100
rect 3500 3900 3900 7100
rect 6800 3900 7200 7100
rect 7500 3900 7900 7100
rect 100 0 500 3200
rect 800 0 1200 3200
rect 2100 0 2500 3200
rect 2800 0 3200 3200
rect 4100 0 4500 3200
rect 4800 0 5200 3200
rect 6100 0 6500 3200
rect 6800 0 7200 3200
rect 7500 0 7900 3200
<< ndiff >>
rect 1700 10900 2000 11000
rect 1700 7900 1800 10900
rect 1900 7900 2000 10900
rect 1700 7800 2000 7900
rect 2400 10900 2700 11000
rect 2400 7900 2500 10900
rect 2600 7900 2700 10900
rect 2400 7800 2700 7900
rect 3100 10900 3400 11000
rect 3100 7900 3200 10900
rect 3300 7900 3400 10900
rect 3100 7800 3400 7900
rect 4600 10900 4900 11000
rect 4600 7900 4700 10900
rect 4800 7900 4900 10900
rect 4600 7800 4900 7900
rect 5300 10900 5600 11000
rect 5300 7900 5400 10900
rect 5500 7900 5600 10900
rect 5300 7800 5600 7900
rect 6000 10900 6300 11000
rect 6000 7900 6100 10900
rect 6200 7900 6300 10900
rect 6000 7800 6300 7900
rect 7200 10900 7500 11000
rect 7200 7900 7300 10900
rect 7400 7900 7500 10900
rect 7200 7800 7500 7900
rect 7900 10900 8200 11000
rect 7900 7900 8000 10900
rect 8100 7900 8200 10900
rect 7900 7800 8200 7900
rect 2500 7000 2800 7100
rect 2500 4000 2600 7000
rect 2700 4000 2800 7000
rect 2500 3900 2800 4000
rect 3200 7000 3500 7100
rect 3200 4000 3300 7000
rect 3400 4000 3500 7000
rect 3200 3900 3500 4000
rect 3900 7000 4200 7100
rect 3900 4000 4000 7000
rect 4100 4000 4200 7000
rect 3900 3900 4200 4000
rect 6500 7000 6800 7100
rect 6500 4000 6600 7000
rect 6700 4000 6800 7000
rect 6500 3900 6800 4000
rect 7200 7000 7500 7100
rect 7200 4000 7300 7000
rect 7400 4000 7500 7000
rect 7200 3900 7500 4000
rect 7900 7000 8200 7100
rect 7900 4000 8000 7000
rect 8100 4000 8200 7000
rect 7900 3900 8200 4000
rect -200 100 -100 3200
rect 0 100 100 3200
rect -200 0 100 100
rect 500 3100 800 3200
rect 500 100 600 3100
rect 700 100 800 3100
rect 500 0 800 100
rect 1200 3100 1500 3200
rect 1800 3100 2100 3200
rect 1200 100 1300 3100
rect 1400 100 1500 3100
rect 1800 100 1900 3100
rect 2000 100 2100 3100
rect 1200 0 1500 100
rect 1800 0 2100 100
rect 2500 3100 2800 3200
rect 2500 100 2600 3100
rect 2700 100 2800 3100
rect 2500 0 2800 100
rect 3200 3100 3500 3200
rect 3800 3100 4100 3200
rect 3200 100 3300 3100
rect 3400 100 3500 3100
rect 3800 100 3900 3100
rect 4000 100 4100 3100
rect 3200 0 3500 100
rect 3800 0 4100 100
rect 4500 3100 4800 3200
rect 4500 100 4600 3100
rect 4700 100 4800 3100
rect 4500 0 4800 100
rect 5200 3100 5500 3200
rect 5800 3100 6100 3200
rect 5200 100 5300 3100
rect 5400 100 5500 3100
rect 5800 100 5900 3100
rect 6000 100 6100 3100
rect 5200 0 5500 100
rect 5800 0 6100 100
rect 6500 3100 6800 3200
rect 6500 100 6600 3100
rect 6700 100 6800 3100
rect 6500 0 6800 100
rect 7200 3100 7500 3200
rect 7200 100 7300 3100
rect 7400 100 7500 3100
rect 7200 0 7500 100
rect 7900 3100 8200 3200
rect 7900 100 8000 3100
rect 8100 100 8200 3100
rect 7900 0 8200 100
<< ndiffc >>
rect 1800 7900 1900 10900
rect 2500 7900 2600 10900
rect 3200 7900 3300 10900
rect 4700 7900 4800 10900
rect 5400 7900 5500 10900
rect 6100 7900 6200 10900
rect 7300 7900 7400 10900
rect 8000 7900 8100 10900
rect 2600 4000 2700 7000
rect 3300 4000 3400 7000
rect 4000 4000 4100 7000
rect 6600 4000 6700 7000
rect 7300 4000 7400 7000
rect 8000 4000 8100 7000
rect -100 100 0 3100
rect 600 100 700 3100
rect 1300 100 1400 3100
rect 1900 100 2000 3100
rect 2600 100 2700 3100
rect 3300 100 3400 3100
rect 3900 100 4000 3100
rect 4600 100 4700 3100
rect 5300 100 5400 3100
rect 5900 100 6000 3100
rect 6600 100 6700 3100
rect 7300 100 7400 3100
rect 8000 100 8100 3100
<< psubdiff >>
rect 1400 10900 1700 11000
rect 1400 7900 1500 10900
rect 1600 7900 1700 10900
rect 1400 7800 1700 7900
rect 3400 10900 3700 11000
rect 3400 7900 3500 10900
rect 3600 7900 3700 10900
rect 3400 7800 3700 7900
rect 4300 10900 4600 11000
rect 4300 7900 4400 10900
rect 4500 7900 4600 10900
rect 4300 7800 4600 7900
rect 6300 10900 6600 11000
rect 6300 7900 6400 10900
rect 6500 7900 6600 10900
rect 6300 7800 6600 7900
rect 8200 10900 8500 11000
rect 8200 7900 8300 10900
rect 8400 7900 8500 10900
rect 8200 7800 8500 7900
rect 2200 7000 2500 7100
rect 2200 4000 2300 7000
rect 2400 4000 2500 7000
rect 2200 3900 2500 4000
rect 4200 7000 4500 7100
rect 4200 4000 4300 7000
rect 4400 4000 4500 7000
rect 4200 3900 4500 4000
rect 6200 7000 6500 7100
rect 6200 4000 6300 7000
rect 6400 4000 6500 7000
rect 6200 3900 6500 4000
rect 8200 7000 8500 7100
rect 8200 4000 8300 7000
rect 8400 4000 8500 7000
rect 8200 3900 8500 4000
rect -500 3100 -200 3200
rect -500 100 -400 3100
rect -300 100 -200 3100
rect -500 0 -200 100
rect 1500 3100 1800 3200
rect 1500 100 1600 3100
rect 1700 100 1800 3100
rect 1500 0 1800 100
rect 3500 3100 3800 3200
rect 3500 100 3600 3100
rect 3700 100 3800 3100
rect 3500 0 3800 100
rect 5500 3100 5800 3200
rect 5500 100 5600 3100
rect 5700 100 5800 3100
rect 5500 0 5800 100
rect 8200 3100 8500 3200
rect 8200 100 8300 3100
rect 8400 100 8500 3100
rect 8200 0 8500 100
<< psubdiffcont >>
rect 1500 7900 1600 10900
rect 3500 7900 3600 10900
rect 4400 7900 4500 10900
rect 6400 7900 6500 10900
rect 8300 7900 8400 10900
rect 2300 4000 2400 7000
rect 4300 4000 4400 7000
rect 6300 4000 6400 7000
rect 8300 4000 8400 7000
rect -400 100 -300 3100
rect 1600 100 1700 3100
rect 3600 100 3700 3100
rect 5600 100 5700 3100
rect 8300 100 8400 3100
<< poly >>
rect 2000 11000 2400 11100
rect 2700 11000 3100 11100
rect 4900 11000 5300 11100
rect 5600 11000 6000 11100
rect 7500 11000 7900 11100
rect 2000 7650 2400 7800
rect 2000 7550 2050 7650
rect 2350 7550 2400 7650
rect 2000 7500 2400 7550
rect 2700 7450 3100 7800
rect 4900 7700 5300 7800
rect 5600 7700 6000 7800
rect 4900 7600 6000 7700
rect 7500 7450 7900 7800
rect 2700 7350 7900 7450
rect 2800 7100 3200 7200
rect 3500 7100 3900 7200
rect 6800 7100 7200 7200
rect 7500 7100 7900 7200
rect 2800 3800 3200 3900
rect 3500 3800 3900 3900
rect 6800 3800 7200 3900
rect 7500 3800 7900 3900
rect 100 3200 500 3300
rect 800 3200 1200 3300
rect 2100 3200 2500 3300
rect 2800 3200 3200 3300
rect 4100 3200 4500 3300
rect 4800 3200 5200 3300
rect 6100 3200 6500 3300
rect 6800 3200 7200 3300
rect 7500 3200 7900 3300
rect 100 -100 500 0
rect 800 -100 1200 0
rect 2100 -100 2500 0
rect 2800 -100 3200 0
rect 4100 -100 4500 0
rect 4800 -100 5200 0
rect 6100 -100 6500 0
rect 6800 -100 7200 0
rect 7500 -100 7900 0
<< polycont >>
rect 2050 7550 2350 7650
<< locali >>
rect 1800 11200 7400 11300
rect 1500 10900 1600 11000
rect 1800 10900 1900 11200
rect 3500 10900 3600 11000
rect 1600 7900 1800 10900
rect 1900 7900 2000 10900
rect 2400 7900 2500 10900
rect 2600 7900 2700 10900
rect 3100 7900 3200 10900
rect 3300 7900 3400 10900
rect 1500 7800 1600 7900
rect 1800 7650 1900 7900
rect 2000 7650 2400 7700
rect 1800 7550 2050 7650
rect 2350 7550 2400 7650
rect 2000 7500 2400 7550
rect 2500 7450 2600 7900
rect 3500 7800 3600 7900
rect 4400 10900 4500 11000
rect 5400 10900 5500 11200
rect 6400 10900 6500 11000
rect 7300 10900 7400 11200
rect 8300 10900 8400 11000
rect 4600 7900 4700 10900
rect 4800 7900 4900 10900
rect 5300 7900 5400 10900
rect 5500 7900 5600 10900
rect 6000 7900 6100 10900
rect 6200 7900 6300 10900
rect 7200 7900 7300 10900
rect 7400 7900 7500 10900
rect 7900 7900 8000 10900
rect 8100 7900 8200 10900
rect 4400 7800 4500 7900
rect 4700 7550 4800 7900
rect 6400 7800 6500 7900
rect 1900 7350 2600 7450
rect 3300 7450 4800 7550
rect 1900 3850 2000 7350
rect 2300 7000 2400 7100
rect 3300 7000 3400 7450
rect 4300 7000 4400 7100
rect 2500 4000 2600 7000
rect 2700 4000 2800 7000
rect 3200 4000 3300 7000
rect 3400 4000 3500 7000
rect 3900 4000 4000 7000
rect 4100 4000 4200 7000
rect 2300 3900 2400 4000
rect 4300 3900 4400 4000
rect 6300 7000 6400 7100
rect 8000 7000 8100 7900
rect 8300 7800 8400 7900
rect 8300 7000 8400 7100
rect 6500 4000 6600 7000
rect 6700 4000 6800 7000
rect 7200 4000 7300 7000
rect 7400 4000 7500 7000
rect 7900 4000 8000 7000
rect 8100 4000 8200 7000
rect 6300 3900 6400 4000
rect 8300 3900 8400 4000
rect -100 3750 2000 3850
rect -400 3100 -300 3200
rect -100 3100 0 3750
rect 1600 3100 1700 3200
rect 3600 3100 3700 3200
rect 5600 3100 5700 3200
rect 8300 3100 8400 3200
rect -200 100 -100 3100
rect 0 100 100 3100
rect 500 100 600 3100
rect 700 100 800 3100
rect 1200 100 1300 3100
rect 1400 100 1500 3100
rect 1800 100 1900 3100
rect 2000 100 2100 3100
rect 2500 100 2600 3100
rect 2700 100 2800 3100
rect 3200 100 3300 3100
rect 3400 100 3500 3100
rect 3800 100 3900 3100
rect 4000 100 4100 3100
rect 4500 100 4600 3100
rect 4700 100 4800 3100
rect 5200 100 5300 3100
rect 5400 100 5500 3100
rect 5800 100 5900 3100
rect 6000 100 6100 3100
rect 6500 100 6600 3100
rect 6700 100 6800 3100
rect 7200 100 7300 3100
rect 7400 100 7500 3100
rect 7900 100 8000 3100
rect 8100 100 8200 3100
rect -400 0 -300 100
rect 1600 0 1700 100
rect 3600 0 3700 100
rect 5600 0 5700 100
rect 8300 0 8400 100
<< viali >>
rect 1500 7900 1600 10900
<< end >>
