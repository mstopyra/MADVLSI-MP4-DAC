magic
tech sky130A
timestamp 1701228941
<< nwell >>
rect -1400 7005 6200 10600
rect -1400 7000 6175 7005
<< nmos >>
rect -1100 3200 -700 6400
rect -400 3200 0 6400
rect 100 3200 500 6400
rect 600 3200 1000 6400
rect 1100 3200 1500 6400
rect 1800 3200 2200 6400
rect 2500 3200 2900 6400
rect 3200 3200 3600 6400
rect 3700 3200 4100 6400
rect 4200 3200 4600 6400
rect 4700 3200 5100 6400
rect 5400 3200 5800 6400
<< pmos >>
rect -1100 7100 -700 10300
rect -375 7100 25 10300
rect 125 7100 525 10300
rect 625 7100 1025 10300
rect 1125 7100 1525 10300
rect 1625 7100 2025 10300
rect 2375 7100 2775 10300
rect 2875 7100 3275 10300
rect 3375 7100 3775 10300
rect 3875 7100 4275 10300
rect 4375 7100 4775 10300
rect 5125 7100 5525 10300
<< ndiff >>
rect -1195 6380 -1100 6400
rect -1195 3220 -1180 6380
rect -1120 3220 -1100 6380
rect -1195 3200 -1100 3220
rect -700 6380 -605 6400
rect -700 3220 -680 6380
rect -620 3220 -605 6380
rect -700 3200 -605 3220
rect -495 6380 -400 6400
rect -495 3220 -480 6380
rect -420 3220 -400 6380
rect -495 3200 -400 3220
rect 0 6380 100 6400
rect 0 3220 20 6380
rect 80 3220 100 6380
rect 0 3200 100 3220
rect 500 6380 600 6400
rect 500 3220 520 6380
rect 580 3220 600 6380
rect 500 3200 600 3220
rect 1000 6380 1100 6400
rect 1000 3220 1020 6380
rect 1080 3220 1100 6380
rect 1000 3200 1100 3220
rect 1500 6380 1595 6400
rect 1500 3220 1520 6380
rect 1580 3220 1595 6380
rect 1500 3200 1595 3220
rect 1705 6380 1800 6400
rect 1705 3220 1720 6380
rect 1780 3220 1800 6380
rect 1705 3200 1800 3220
rect 2200 6380 2500 6400
rect 2200 3220 2220 6380
rect 2480 3220 2500 6380
rect 2200 3200 2500 3220
rect 2900 6380 2995 6400
rect 2900 3220 2920 6380
rect 2980 3220 2995 6380
rect 2900 3200 2995 3220
rect 3105 6380 3200 6400
rect 3105 3220 3120 6380
rect 3180 3220 3200 6380
rect 3105 3200 3200 3220
rect 3600 6380 3700 6400
rect 3600 3220 3620 6380
rect 3680 3220 3700 6380
rect 3600 3200 3700 3220
rect 4100 6380 4200 6400
rect 4100 3220 4120 6380
rect 4180 3220 4200 6380
rect 4100 3200 4200 3220
rect 4600 6380 4700 6400
rect 4600 3220 4620 6380
rect 4680 3220 4700 6380
rect 4600 3200 4700 3220
rect 5100 6380 5195 6400
rect 5100 3220 5120 6380
rect 5180 3220 5195 6380
rect 5100 3200 5195 3220
rect 5305 6380 5400 6400
rect 5305 3220 5320 6380
rect 5380 3220 5400 6380
rect 5305 3200 5400 3220
rect 5800 6380 5895 6400
rect 5800 3220 5820 6380
rect 5880 3220 5895 6380
rect 5800 3200 5895 3220
<< pdiff >>
rect -1200 10280 -1100 10300
rect -1200 7120 -1180 10280
rect -1120 7120 -1100 10280
rect -1200 7100 -1100 7120
rect -700 10280 -600 10300
rect -700 7120 -680 10280
rect -620 7120 -600 10280
rect -700 7100 -600 7120
rect -475 10280 -375 10300
rect -475 7120 -455 10280
rect -395 7120 -375 10280
rect -475 7100 -375 7120
rect 25 7100 125 10300
rect 525 7100 625 10300
rect 1025 7100 1125 10300
rect 1525 7100 1625 10300
rect 2025 10280 2125 10300
rect 2025 7120 2045 10280
rect 2105 7120 2125 10280
rect 2025 7100 2125 7120
rect 2280 10280 2375 10300
rect 2280 7120 2295 10280
rect 2355 7120 2375 10280
rect 2280 7100 2375 7120
rect 2775 7100 2875 10300
rect 3275 7100 3375 10300
rect 3775 7100 3875 10300
rect 4275 7100 4375 10300
rect 4775 10280 4875 10300
rect 4775 7120 4795 10280
rect 4855 7120 4875 10280
rect 4775 7100 4875 7120
rect 5030 10280 5125 10300
rect 5030 7120 5045 10280
rect 5105 7120 5125 10280
rect 5030 7100 5125 7120
rect 5525 10280 5625 10300
rect 5525 7120 5545 10280
rect 5605 7120 5625 10280
rect 5525 7100 5625 7120
<< ndiffc >>
rect -1180 3220 -1120 6380
rect -680 3220 -620 6380
rect -480 3220 -420 6380
rect 20 3220 80 6380
rect 520 3220 580 6380
rect 1020 3220 1080 6380
rect 1520 3220 1580 6380
rect 1720 3220 1780 6380
rect 2220 3220 2480 6380
rect 2920 3220 2980 6380
rect 3120 3220 3180 6380
rect 3620 3220 3680 6380
rect 4120 3220 4180 6380
rect 4620 3220 4680 6380
rect 5120 3220 5180 6380
rect 5320 3220 5380 6380
rect 5820 3220 5880 6380
<< pdiffc >>
rect -1180 7120 -1120 10280
rect -680 7120 -620 10280
rect -455 7120 -395 10280
rect 2045 7120 2105 10280
rect 2295 7120 2355 10280
rect 4795 7120 4855 10280
rect 5045 7120 5105 10280
rect 5545 7120 5605 10280
<< psubdiff >>
rect -1275 6390 -1225 6395
rect -1275 3215 -1260 6390
rect -1240 3215 -1225 6390
rect -1275 3200 -1225 3215
rect -575 6390 -525 6395
rect -575 3215 -560 6390
rect -540 3215 -525 6390
rect -575 3200 -525 3215
rect 1625 6390 1675 6395
rect 1625 3215 1640 6390
rect 1660 3215 1675 6390
rect 1625 3200 1675 3215
rect 3025 6390 3075 6395
rect 3025 3215 3040 6390
rect 3060 3215 3075 6390
rect 3025 3200 3075 3215
rect 5225 6390 5275 6395
rect 5225 3215 5240 6390
rect 5260 3215 5275 6390
rect 5225 3200 5275 3215
rect 5925 6390 5975 6395
rect 5925 3215 5940 6390
rect 5960 3215 5975 6390
rect 5925 3200 5975 3215
<< nsubdiff >>
rect -570 10290 -505 10300
rect -570 7115 -555 10290
rect -520 7115 -505 10290
rect -570 7100 -505 7115
rect 2155 10280 2250 10300
rect 2155 7120 2170 10280
rect 2230 7120 2250 10280
rect 2155 7100 2250 7120
rect 4905 10280 5000 10300
rect 4905 7120 4920 10280
rect 4980 7120 5000 10280
rect 4905 7100 5000 7120
<< psubdiffcont >>
rect -1260 3215 -1240 6390
rect -560 3215 -540 6390
rect 1640 3215 1660 6390
rect 3040 3215 3060 6390
rect 5240 3215 5260 6390
rect 5940 3215 5960 6390
<< nsubdiffcont >>
rect -555 7115 -520 10290
rect 2170 7120 2230 10280
rect 4920 7120 4980 10280
<< poly >>
rect -1400 10400 5425 10500
rect -1000 10325 -800 10400
rect -275 10325 -75 10400
rect 225 10325 425 10400
rect 725 10325 925 10400
rect 1225 10325 1425 10400
rect 1725 10325 1925 10400
rect 2475 10325 2675 10400
rect 2975 10325 3175 10400
rect 3475 10325 3675 10400
rect 3975 10325 4175 10400
rect 4475 10325 4675 10400
rect 5225 10325 5425 10400
rect -1100 10300 -700 10325
rect -375 10300 25 10325
rect 125 10300 525 10325
rect 625 10300 1025 10325
rect 1125 10300 1525 10325
rect 1625 10300 2025 10325
rect 2375 10300 2775 10325
rect 2875 10300 3275 10325
rect 3375 10300 3775 10325
rect 3875 10300 4275 10325
rect 4375 10300 4775 10325
rect 5125 10300 5525 10325
rect -1100 7075 -700 7100
rect -375 7075 25 7100
rect 125 7075 525 7100
rect 625 7075 1025 7100
rect 1125 7075 1525 7100
rect 1625 7075 2025 7100
rect 2375 7075 2775 7100
rect 2875 7075 3275 7100
rect 3375 7075 3775 7100
rect 3875 7075 4275 7100
rect 4375 7075 4775 7100
rect 5125 7075 5525 7100
rect 2000 6980 2200 7000
rect 2000 6920 2120 6980
rect 2180 6920 2200 6980
rect 2000 6900 2200 6920
rect 2000 6700 2100 6900
rect -1200 6590 -1000 6600
rect -1200 6510 -1190 6590
rect -1110 6510 -1000 6590
rect -1200 6500 -1000 6510
rect -1100 6420 -1000 6500
rect 1200 6500 3500 6700
rect 1200 6420 1400 6500
rect 1900 6420 2100 6500
rect 2600 6420 2800 6500
rect 3300 6420 3500 6500
rect 5700 6590 5900 6600
rect 5700 6510 5810 6590
rect 5890 6510 5900 6590
rect 5700 6500 5900 6510
rect 5700 6420 5800 6500
rect -1100 6400 -700 6420
rect -400 6400 0 6420
rect 100 6400 500 6420
rect 600 6400 1000 6420
rect 1100 6400 1500 6420
rect 1800 6400 2200 6420
rect 2500 6400 2900 6420
rect 3200 6400 3600 6420
rect 3700 6400 4100 6420
rect 4200 6400 4600 6420
rect 4700 6400 5100 6420
rect 5400 6400 5800 6420
rect -1100 3180 -700 3200
rect -400 3180 0 3200
rect 100 3180 500 3200
rect 600 3180 1000 3200
rect 1100 3180 1500 3200
rect 1800 3180 2200 3200
rect 2500 3180 2900 3200
rect 3200 3180 3600 3200
rect 3700 3180 4100 3200
rect 4200 3180 4600 3200
rect 4700 3180 5100 3200
rect 5400 3180 5800 3200
rect -200 3050 0 3180
rect -200 2950 -150 3050
rect -50 2950 0 3050
rect -200 2900 0 2950
rect 200 3050 400 3180
rect 200 2950 250 3050
rect 350 2950 400 3050
rect 200 2900 400 2950
rect 700 3050 900 3180
rect 700 2950 750 3050
rect 850 2950 900 3050
rect 700 2900 900 2950
rect 1100 3050 1300 3180
rect 1100 2950 1150 3050
rect 1250 2950 1300 3050
rect 1100 2900 1300 2950
rect 3400 3050 3600 3180
rect 3400 2950 3450 3050
rect 3550 2950 3600 3050
rect 3400 2900 3600 2950
rect 3800 3050 4000 3180
rect 3800 2950 3850 3050
rect 3950 2950 4000 3050
rect 3800 2900 4000 2950
rect 4300 3050 4500 3180
rect 4300 2950 4350 3050
rect 4450 2950 4500 3050
rect 4300 2900 4500 2950
rect 4700 3050 4900 3180
rect 4700 2950 4750 3050
rect 4850 2950 4900 3050
rect 4700 2900 4900 2950
<< polycont >>
rect 2120 6920 2180 6980
rect -1190 6510 -1110 6590
rect 5810 6510 5890 6590
rect -150 2950 -50 3050
rect 250 2950 350 3050
rect 750 2950 850 3050
rect 1150 2950 1250 3050
rect 3450 2950 3550 3050
rect 3850 2950 3950 3050
rect 4350 2950 4450 3050
rect 4750 2950 4850 3050
<< locali >>
rect -1190 10280 -1110 10300
rect -1190 7120 -1180 10280
rect -1120 7120 -1110 10280
rect -1190 7000 -1110 7120
rect -690 10280 -610 10300
rect -690 7120 -680 10280
rect -620 7120 -610 10280
rect -690 7100 -610 7120
rect -570 10290 -505 10300
rect -570 7115 -555 10290
rect -520 7115 -505 10290
rect -570 7100 -505 7115
rect -465 10280 -385 10300
rect -465 7120 -455 10280
rect -395 7120 -385 10280
rect -465 7110 -385 7120
rect 2035 10280 2115 10300
rect 2035 7120 2045 10280
rect 2105 7120 2115 10280
rect 2035 7080 2115 7120
rect 2160 10280 2240 10300
rect 2160 7120 2170 10280
rect 2230 7120 2240 10280
rect 2160 7100 2240 7120
rect 2285 10280 2365 10300
rect 2285 7120 2295 10280
rect 2355 7120 2365 10280
rect 2285 7080 2365 7120
rect 4785 10290 4865 10300
rect 5035 10290 5115 10300
rect 4785 10280 4875 10290
rect 4785 7120 4795 10280
rect 4855 7120 4875 10280
rect 4785 7110 4875 7120
rect 4905 10280 5000 10290
rect 4905 7120 4920 10280
rect 4980 7120 5000 10280
rect 4905 7110 5000 7120
rect 5030 10280 5115 10290
rect 5030 7120 5045 10280
rect 5105 7120 5115 10280
rect 5030 7110 5115 7120
rect 5535 10280 5615 10300
rect 5535 7120 5545 10280
rect 5605 7120 5615 10280
rect 2035 7000 2365 7080
rect 5535 7000 5615 7120
rect -1200 6800 -1100 7000
rect 2100 6980 2200 7000
rect 2100 6920 2120 6980
rect 2180 6920 2200 6980
rect 2100 6900 2200 6920
rect 5525 6800 5625 7000
rect -1400 6700 5900 6800
rect -1200 6590 -1100 6700
rect -1200 6510 -1190 6590
rect -1110 6510 -1100 6590
rect -1200 6500 -1100 6510
rect -700 6500 5400 6600
rect 5800 6590 5900 6700
rect 5800 6510 5810 6590
rect 5890 6510 5900 6590
rect 5800 6500 5900 6510
rect -1270 3215 -1260 6390
rect -1240 3215 -1230 6390
rect -1270 3205 -1230 3215
rect -1190 6380 -1110 6500
rect -1190 3220 -1180 6380
rect -1120 3220 -1110 6380
rect -1190 3210 -1110 3220
rect -690 6380 -610 6500
rect -690 3220 -680 6380
rect -620 3220 -610 6380
rect -690 3210 -610 3220
rect -570 3215 -560 6390
rect -540 3215 -530 6390
rect -570 3205 -530 3215
rect -490 6380 -410 6500
rect -490 3220 -480 6380
rect -420 3220 -410 6380
rect -490 3210 -410 3220
rect 10 6380 90 6390
rect 10 3220 20 6380
rect 80 3220 90 6380
rect 10 3100 90 3220
rect 510 6380 590 6390
rect 510 3220 520 6380
rect 580 3220 590 6380
rect 510 3100 590 3220
rect 1010 6380 1090 6390
rect 1010 3220 1020 6380
rect 1080 3220 1090 6380
rect 1010 3100 1090 3220
rect 1510 6380 1590 6500
rect 1510 3220 1520 6380
rect 1580 3220 1590 6380
rect 1510 3210 1590 3220
rect 1630 3215 1640 6390
rect 1660 3215 1670 6390
rect 1630 3205 1670 3215
rect 1710 6380 1790 6500
rect 1710 3220 1720 6380
rect 1780 3220 1790 6380
rect 1710 3210 1790 3220
rect 2200 6380 2500 6400
rect 2200 3220 2220 6380
rect 2480 3220 2500 6380
rect 2200 3200 2500 3220
rect 2910 6380 2990 6500
rect 2910 3220 2920 6380
rect 2980 3220 2990 6380
rect 2910 3210 2990 3220
rect 3030 3215 3040 6390
rect 3060 3215 3070 6390
rect 3030 3205 3070 3215
rect 3110 6380 3190 6500
rect 3110 3220 3120 6380
rect 3180 3220 3190 6380
rect 3110 3210 3190 3220
rect 3610 6380 3690 6390
rect 3610 3220 3620 6380
rect 3680 3220 3690 6380
rect 3610 3100 3690 3220
rect 4110 6380 4190 6390
rect 4110 3220 4120 6380
rect 4180 3220 4190 6380
rect 4110 3100 4190 3220
rect 4610 6380 4690 6390
rect 4610 3220 4620 6380
rect 4680 3220 4690 6380
rect 4610 3100 4690 3220
rect 5110 6380 5190 6500
rect 5110 3220 5120 6380
rect 5180 3220 5190 6380
rect 5110 3210 5190 3220
rect 5230 3215 5240 6390
rect 5260 3215 5270 6390
rect 5230 3205 5270 3215
rect 5310 6380 5390 6500
rect 5310 3220 5320 6380
rect 5380 3220 5390 6380
rect 5310 3210 5390 3220
rect 5810 6380 5890 6500
rect 5810 3220 5820 6380
rect 5880 3220 5890 6380
rect 5810 3210 5890 3220
rect 5930 3215 5940 6390
rect 5960 3215 5970 6390
rect 5930 3205 5970 3215
rect -200 3050 1300 3100
rect -200 2950 -150 3050
rect -50 2950 250 3050
rect 350 2950 750 3050
rect 850 2950 1150 3050
rect 1250 2950 1300 3050
rect -200 2900 1300 2950
rect 3400 3050 4900 3100
rect 3400 2950 3450 3050
rect 3550 2950 3850 3050
rect 3950 2950 4350 3050
rect 4450 2950 4750 3050
rect 4850 2950 4900 3050
rect 3400 2900 4900 2950
<< viali >>
rect -555 7115 -520 10290
rect 2170 7120 2230 10280
rect 4920 7120 4980 10280
rect -1260 3215 -1240 6390
rect -560 3215 -540 6390
rect 1640 3215 1660 6390
rect 2220 3220 2480 6380
rect 3040 3215 3060 6390
rect 5240 3215 5260 6390
rect 5940 3215 5960 6390
<< metal1 >>
rect 2125 10300 2155 10305
rect 2250 10300 2280 10305
rect -1400 10290 6200 10300
rect -1400 7115 -555 10290
rect -520 10280 6200 10290
rect -520 7120 2170 10280
rect 2230 7120 4920 10280
rect 4980 7120 6200 10280
rect -520 7115 6200 7120
rect -1400 7100 6200 7115
rect -1400 6390 6100 6400
rect -1400 3215 -1260 6390
rect -1240 3215 -560 6390
rect -540 3215 1640 6390
rect 1660 6380 3040 6390
rect 1660 3220 2220 6380
rect 2480 3220 3040 6380
rect 1660 3215 3040 3220
rect 3060 3215 5240 6390
rect 5260 3215 5940 6390
rect 5960 3215 6100 6390
rect -1400 3200 6100 3215
<< labels >>
flabel metal1 -1400 8600 -1395 8605 0 FreeSans 800 0 0 0 VP
port 1 nsew
flabel metal1 -1400 4600 -1395 4605 0 FreeSans 800 0 0 0 VN
port 2 nsew
flabel poly -1400 10450 -1400 10450 0 FreeSans 800 0 0 0 VBP
port 3 nsew
flabel locali -1400 6750 -1400 6750 0 FreeSans 800 0 0 0 VCN
port 4 nsew
<< end >>
