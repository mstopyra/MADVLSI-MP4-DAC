magic
tech sky130A
timestamp 1701115757
<< nwell >>
rect -1400 -800 6500 7200
<< pmos >>
rect -500 3400 -100 6600
rect 1200 3400 1600 6600
rect 1900 3400 2300 6600
rect 3300 3400 3700 6600
rect -500 -200 -100 3000
rect 1200 -200 1600 3000
rect 1900 -200 2300 3000
rect 3300 -200 3700 3000
<< pdiff >>
rect -800 6500 -500 6600
rect -800 3500 -700 6500
rect -600 3500 -500 6500
rect -800 3400 -500 3500
rect -100 6500 200 6600
rect -100 3500 0 6500
rect 100 3500 200 6500
rect -100 3400 200 3500
rect 900 6500 1200 6600
rect 900 3500 1000 6500
rect 1100 3500 1200 6500
rect 900 3400 1200 3500
rect 1600 6500 1900 6600
rect 1600 3500 1700 6500
rect 1800 3500 1900 6500
rect 1600 3400 1900 3500
rect 2300 6500 2600 6600
rect 3000 6500 3300 6600
rect 2300 3500 2400 6500
rect 2500 3500 2600 6500
rect 3000 3500 3100 6500
rect 3200 3500 3300 6500
rect 2300 3400 2600 3500
rect 3000 3400 3300 3500
rect 3700 6500 4000 6600
rect 3700 3500 3800 6500
rect 3900 3500 4000 6500
rect 3700 3400 4000 3500
rect -800 2900 -500 3000
rect -800 -100 -700 2900
rect -600 -100 -500 2900
rect -800 -200 -500 -100
rect -100 2900 200 3000
rect -100 -100 0 2900
rect 100 -100 200 2900
rect -100 -200 200 -100
rect 900 2900 1200 3000
rect 900 -100 1000 2900
rect 1100 -100 1200 2900
rect 900 -200 1200 -100
rect 1600 2900 1900 3000
rect 1600 -100 1700 2900
rect 1800 -100 1900 2900
rect 1600 -200 1900 -100
rect 2300 2900 2600 3000
rect 3000 2900 3300 3000
rect 2300 -100 2400 2900
rect 2500 -100 2600 2900
rect 3000 -100 3100 2900
rect 3200 -100 3300 2900
rect 2300 -200 2600 -100
rect 3000 -200 3300 -100
rect 3700 2900 4000 3000
rect 3700 -100 3800 2900
rect 3900 -100 4000 2900
rect 3700 -200 4000 -100
<< pdiffc >>
rect -700 3500 -600 6500
rect 0 3500 100 6500
rect 1000 3500 1100 6500
rect 1700 3500 1800 6500
rect 2400 3500 2500 6500
rect 3100 3500 3200 6500
rect 3800 3500 3900 6500
rect -700 -100 -600 2900
rect 0 -100 100 2900
rect 1000 -100 1100 2900
rect 1700 -100 1800 2900
rect 2400 -100 2500 2900
rect 3100 -100 3200 2900
rect 3800 -100 3900 2900
<< nsubdiff >>
rect -1200 6500 -800 6600
rect -1200 3500 -1100 6500
rect -900 3500 -800 6500
rect -1200 3400 -800 3500
rect 500 6500 900 6600
rect 500 3500 600 6500
rect 800 3500 900 6500
rect 500 3400 900 3500
rect 2600 6500 3000 6600
rect 2600 3500 2700 6500
rect 2900 3500 3000 6500
rect 2600 3400 3000 3500
rect -1200 2900 -800 3000
rect -1200 -100 -1100 2900
rect -900 -100 -800 2900
rect -1200 -200 -800 -100
rect 500 2900 900 3000
rect 500 -100 600 2900
rect 800 -100 900 2900
rect 500 -200 900 -100
rect 2600 2900 3000 3000
rect 2600 -100 2700 2900
rect 2900 -100 3000 2900
rect 2600 -200 3000 -100
<< nsubdiffcont >>
rect -1100 3500 -900 6500
rect 600 3500 800 6500
rect 2700 3500 2900 6500
rect -1100 -100 -900 2900
rect 600 -100 800 2900
rect 2700 -100 2900 2900
<< poly >>
rect 3300 6850 3700 6900
rect -500 6750 -100 6800
rect -500 6650 -450 6750
rect -150 6650 -100 6750
rect -500 6600 -100 6650
rect 1200 6750 1600 6800
rect 1200 6650 1250 6750
rect 1550 6650 1600 6750
rect 1200 6600 1600 6650
rect 1900 6750 2300 6800
rect 1900 6650 1950 6750
rect 2250 6650 2300 6750
rect 1900 6600 2300 6650
rect 3300 6750 3350 6850
rect 3650 6750 3700 6850
rect 3300 6600 3700 6750
rect -500 3300 -100 3400
rect -500 3150 -100 3200
rect -500 3050 -450 3150
rect -150 3050 -100 3150
rect -500 3000 -100 3050
rect 1200 3000 1600 3400
rect 1900 3000 2300 3400
rect 3300 3350 3700 3400
rect 3300 3250 3700 3300
rect 3300 3150 3350 3250
rect 3650 3150 3700 3250
rect 3300 3000 3700 3150
rect -500 -300 -100 -200
rect 1200 -300 1600 -200
rect 1900 -300 2300 -200
rect 3300 -300 3700 -200
<< polycont >>
rect -450 6650 -150 6750
rect 1250 6650 1550 6750
rect 1950 6650 2250 6750
rect 3350 6750 3650 6850
rect -450 3050 -150 3150
rect 3350 3150 3650 3250
<< locali >>
rect 3000 6800 3200 6900
rect -800 6750 -100 6800
rect -800 6650 -450 6750
rect -150 6650 -100 6750
rect -800 6600 -100 6650
rect 1200 6750 1600 6800
rect 1200 6650 1250 6750
rect 1550 6700 1600 6750
rect 1900 6750 2300 6800
rect 1900 6700 1950 6750
rect 1550 6650 1950 6700
rect 2250 6650 2300 6750
rect 1200 6600 2300 6650
rect -1100 6500 -600 6600
rect -1200 3500 -1100 3600
rect -900 3500 -700 6500
rect -1200 3400 -600 3500
rect 0 6500 100 6600
rect 500 6500 900 6600
rect 500 6400 600 6500
rect 0 3200 100 3500
rect 500 3500 600 3600
rect 800 6400 900 6500
rect 1000 6500 1100 6600
rect 800 3500 900 3600
rect 500 3400 900 3500
rect 1000 3200 1100 3500
rect 1700 6500 1800 6600
rect 1700 3400 1800 3500
rect 2400 6500 2500 6600
rect 2600 6500 3000 6600
rect 2600 6400 2700 6500
rect -800 3150 -100 3200
rect -800 3050 -450 3150
rect -150 3050 -100 3150
rect -800 3000 -100 3050
rect 0 3100 1100 3200
rect -1100 2900 -600 3000
rect -1200 -100 -1100 0
rect -900 -100 -700 2900
rect -1200 -200 -600 -100
rect 0 -200 100 3100
rect 500 2900 900 3000
rect 500 2800 600 2900
rect 500 -100 600 0
rect 800 2800 900 2900
rect 1000 2900 1100 3100
rect 1600 3350 1900 3400
rect 1600 3050 1650 3350
rect 1850 3050 1900 3350
rect 1600 3000 1900 3050
rect 2400 3300 2500 3500
rect 2600 3500 2700 3600
rect 2900 6400 3000 6500
rect 3100 6500 3200 6800
rect 3300 6850 3700 6900
rect 3300 6750 3350 6850
rect 3650 6750 3700 6850
rect 3300 6700 3700 6750
rect 2900 3500 3000 3600
rect 2600 3400 3000 3500
rect 3100 3400 3200 3500
rect 3750 6500 3950 6550
rect 3750 3500 3800 6500
rect 3900 3500 3950 6500
rect 3750 3450 3950 3500
rect 2400 3200 3200 3300
rect 800 -100 900 0
rect 500 -200 900 -100
rect 1000 -300 1100 -100
rect 1700 2900 1800 3000
rect 1700 -200 1800 -100
rect 2400 2900 2500 3200
rect 2600 2900 3000 3000
rect 2600 2800 2700 2900
rect 2400 -300 2500 -100
rect 2600 -100 2700 0
rect 2900 2800 3000 2900
rect 3100 2900 3200 3200
rect 3300 3250 3700 3300
rect 3300 3150 3350 3250
rect 3650 3150 3700 3250
rect 3300 3100 3700 3150
rect 2900 -100 3000 0
rect 2600 -200 3000 -100
rect 3100 -300 3200 -100
rect 3750 2900 3950 2950
rect 3750 -100 3800 2900
rect 3900 -100 3950 2900
rect 3750 -150 3950 -100
rect 1000 -400 2500 -300
<< viali >>
rect -1100 3500 -900 6500
rect 600 3500 800 6500
rect -1100 -100 -900 2900
rect 600 -100 800 2900
rect 1650 3050 1850 3350
rect 2700 3500 2900 6500
rect 2700 -100 2900 2900
rect 3350 3150 3650 3250
rect 3800 -100 3900 2900
<< metal1 >>
rect -1150 6500 -850 6550
rect -1150 3500 -1100 6500
rect -900 3500 -850 6500
rect -1150 3450 -850 3500
rect 550 6500 850 6550
rect 550 3500 600 6500
rect 800 3500 850 6500
rect 550 3450 850 3500
rect 2650 6500 2950 6550
rect 2650 3500 2700 6500
rect 2900 3500 2950 6500
rect 2650 3450 2950 3500
rect 1600 3350 1900 3400
rect 1600 3050 1650 3350
rect 1850 3300 1900 3350
rect 1850 3250 3700 3300
rect 1850 3150 3350 3250
rect 3650 3150 3700 3250
rect 1850 3100 3700 3150
rect 1850 3050 1900 3100
rect 1600 3000 1900 3050
rect -1150 2900 -850 2950
rect -1150 -100 -1100 2900
rect -900 -100 -850 2900
rect -1150 -150 -850 -100
rect 550 2900 850 2950
rect 550 -100 600 2900
rect 800 -100 850 2900
rect 550 -150 850 -100
rect 2650 2900 2950 2950
rect 2650 -100 2700 2900
rect 2900 -100 2950 2900
rect 2650 -150 2950 -100
rect 3750 2900 3950 2950
rect 3750 -100 3800 2900
rect 3900 -100 3950 2900
rect 3750 -150 3950 -100
<< via1 >>
rect -1100 3500 -900 6500
rect 600 3500 800 6500
rect 2700 3500 2900 6500
rect -1100 -100 -900 2900
rect 600 -100 800 2900
rect 2700 -100 2900 2900
rect 3800 -100 3900 2900
<< metal2 >>
rect -1150 6500 -850 6550
rect -1150 3500 -1100 6500
rect -900 3500 -850 6500
rect -1150 2900 -850 3500
rect -1150 -100 -1100 2900
rect -900 -100 -850 2900
rect -1150 -150 -850 -100
rect 550 6500 850 6550
rect 550 3500 600 6500
rect 800 3500 850 6500
rect 550 2900 850 3500
rect 550 -100 600 2900
rect 800 -100 850 2900
rect 550 -150 850 -100
rect 2650 6500 2950 6550
rect 2650 3500 2700 6500
rect 2900 3500 2950 6500
rect 2650 2900 2950 3500
rect 2650 -100 2700 2900
rect 2900 -100 2950 2900
rect 2650 -150 2950 -100
rect 3750 2900 3950 2950
rect 3750 -100 3800 2900
rect 3900 -100 3950 2900
rect 3750 -150 3950 -100
rect -1150 -350 3950 -150
<< end >>
