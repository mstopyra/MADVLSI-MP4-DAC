magic
tech sky130A
timestamp 1700966227
<< nwell >>
rect -8900 -200 21400 4200
<< nmos >>
rect -7200 -5000 -6800 -1800
rect -5800 -5000 -5400 -1800
rect -4400 -5000 -4000 -1800
rect -900 -5000 -500 -1800
rect 500 -5000 900 -1800
rect 4000 -5000 4400 -1800
rect 4500 -5000 4900 -1800
rect 7500 -5000 7900 -1800
rect 8000 -5000 8400 -1800
rect 11500 -5000 11900 -1800
rect 12900 -5000 13300 -1800
rect 16400 -5000 16800 -1800
rect 17800 -5000 18200 -1800
rect 19200 -5000 19600 -1800
<< pmos >>
rect -5200 400 -4800 3600
rect -3800 400 -3400 3600
rect -3300 400 -2900 3600
rect 200 400 600 3600
rect 700 400 1100 3600
rect 4100 400 4500 3600
rect 4600 400 5000 3600
rect 7400 400 7800 3600
rect 7900 400 8300 3600
rect 11300 400 11700 3600
rect 11800 400 12200 3600
rect 15300 400 15700 3600
rect 15800 400 16200 3600
rect 17200 400 17600 3600
<< ndiff >>
rect -8100 -1900 -7200 -1800
rect -8100 -4900 -8000 -1900
rect -7400 -4900 -7200 -1900
rect -8100 -5000 -7200 -4900
rect -6800 -1900 -5800 -1800
rect -6800 -4900 -6600 -1900
rect -6000 -4900 -5800 -1900
rect -6800 -5000 -5800 -4900
rect -5400 -1900 -4400 -1800
rect -5400 -4900 -5200 -1900
rect -4600 -4900 -4400 -1900
rect -5400 -5000 -4400 -4900
rect -4000 -1900 -3100 -1800
rect -4000 -4900 -3800 -1900
rect -3200 -4900 -3100 -1900
rect -4000 -5000 -3100 -4900
rect -1800 -1900 -900 -1800
rect -1800 -4900 -1700 -1900
rect -1100 -4900 -900 -1900
rect -1800 -5000 -900 -4900
rect -500 -1900 500 -1800
rect -500 -4900 -300 -1900
rect 300 -4900 500 -1900
rect -500 -5000 500 -4900
rect 900 -1900 1800 -1800
rect 900 -4900 1100 -1900
rect 1700 -4900 1800 -1900
rect 900 -5000 1800 -4900
rect 3100 -1900 4000 -1800
rect 3100 -4900 3200 -1900
rect 3800 -4900 4000 -1900
rect 3100 -5000 4000 -4900
rect 4400 -5000 4500 -1800
rect 4900 -1900 5900 -1800
rect 4900 -4900 5100 -1900
rect 5700 -4900 5900 -1900
rect 4900 -5000 5900 -4900
rect 6500 -1900 7500 -1800
rect 6500 -4900 6700 -1900
rect 7300 -4900 7500 -1900
rect 6500 -5000 7500 -4900
rect 7900 -5000 8000 -1800
rect 8400 -1900 9300 -1800
rect 8400 -4900 8600 -1900
rect 9200 -4900 9300 -1900
rect 8400 -5000 9300 -4900
rect 10600 -1900 11500 -1800
rect 10600 -4900 10700 -1900
rect 11300 -4900 11500 -1900
rect 10600 -5000 11500 -4900
rect 11900 -1900 12900 -1800
rect 11900 -4900 12100 -1900
rect 12700 -4900 12900 -1900
rect 11900 -5000 12900 -4900
rect 13300 -1900 14200 -1800
rect 13300 -4900 13500 -1900
rect 14100 -4900 14200 -1900
rect 13300 -5000 14200 -4900
rect 15500 -1900 16400 -1800
rect 15500 -4900 15600 -1900
rect 16200 -4900 16400 -1900
rect 15500 -5000 16400 -4900
rect 16800 -1900 17800 -1800
rect 16800 -4900 17000 -1900
rect 17600 -4900 17800 -1900
rect 16800 -5000 17800 -4900
rect 18200 -1900 19200 -1800
rect 18200 -4900 18400 -1900
rect 19000 -4900 19200 -1900
rect 18200 -5000 19200 -4900
rect 19600 -1900 20500 -1800
rect 19600 -4900 19800 -1900
rect 20400 -4900 20500 -1900
rect 19600 -5000 20500 -4900
<< pdiff >>
rect -6100 3500 -5200 3600
rect -6100 500 -6000 3500
rect -5400 500 -5200 3500
rect -6100 400 -5200 500
rect -4800 3500 -3800 3600
rect -4800 500 -4600 3500
rect -4000 500 -3800 3500
rect -4800 400 -3800 500
rect -3400 400 -3300 3600
rect -2900 3500 -2000 3600
rect -2900 500 -2700 3500
rect -2100 500 -2000 3500
rect -2900 400 -2000 500
rect -700 3500 200 3600
rect -700 500 -600 3500
rect 0 500 200 3500
rect -700 400 200 500
rect 600 400 700 3600
rect 1100 3500 2000 3600
rect 1100 500 1300 3500
rect 1900 500 2000 3500
rect 1100 400 2000 500
rect 3200 3500 4100 3600
rect 3200 500 3300 3500
rect 3900 500 4100 3500
rect 3200 400 4100 500
rect 4500 400 4600 3600
rect 5000 3500 5900 3600
rect 5000 500 5200 3500
rect 5800 500 5900 3500
rect 5000 400 5900 500
rect 6500 3500 7400 3600
rect 6500 500 6600 3500
rect 7200 500 7400 3500
rect 6500 400 7400 500
rect 7800 400 7900 3600
rect 8300 3500 9200 3600
rect 8300 500 8500 3500
rect 9100 500 9200 3500
rect 8300 400 9200 500
rect 10400 3500 11300 3600
rect 10400 500 10500 3500
rect 11100 500 11300 3500
rect 10400 400 11300 500
rect 11700 400 11800 3600
rect 12200 3500 13100 3600
rect 12200 500 12400 3500
rect 13000 500 13100 3500
rect 12200 400 13100 500
rect 14400 3500 15300 3600
rect 14400 500 14500 3500
rect 15100 500 15300 3500
rect 14400 400 15300 500
rect 15700 400 15800 3600
rect 16200 3500 17200 3600
rect 16200 500 16400 3500
rect 17000 500 17200 3500
rect 16200 400 17200 500
rect 17600 3500 18500 3600
rect 17600 500 17800 3500
rect 18400 500 18500 3500
rect 17600 400 18500 500
<< ndiffc >>
rect -8000 -4900 -7400 -1900
rect -6600 -4900 -6000 -1900
rect -5200 -4900 -4600 -1900
rect -3800 -4900 -3200 -1900
rect -1700 -4900 -1100 -1900
rect -300 -4900 300 -1900
rect 1100 -4900 1700 -1900
rect 3200 -4900 3800 -1900
rect 5100 -4900 5700 -1900
rect 6700 -4900 7300 -1900
rect 8600 -4900 9200 -1900
rect 10700 -4900 11300 -1900
rect 12100 -4900 12700 -1900
rect 13500 -4900 14100 -1900
rect 15600 -4900 16200 -1900
rect 17000 -4900 17600 -1900
rect 18400 -4900 19000 -1900
rect 19800 -4900 20400 -1900
<< pdiffc >>
rect -6000 500 -5400 3500
rect -4600 500 -4000 3500
rect -2700 500 -2100 3500
rect -600 500 0 3500
rect 1300 500 1900 3500
rect 3300 500 3900 3500
rect 5200 500 5800 3500
rect 6600 500 7200 3500
rect 8500 500 9100 3500
rect 10500 500 11100 3500
rect 12400 500 13000 3500
rect 14500 500 15100 3500
rect 16400 500 17000 3500
rect 17800 500 18400 3500
<< psubdiff >>
rect -8900 -1900 -8100 -1800
rect -8900 -4900 -8800 -1900
rect -8200 -4900 -8100 -1900
rect -8900 -5000 -8100 -4900
rect -2600 -1900 -1800 -1800
rect -2600 -4900 -2500 -1900
rect -1900 -4900 -1800 -1900
rect -2600 -5000 -1800 -4900
rect 2300 -1900 3100 -1800
rect 2300 -4900 2400 -1900
rect 3000 -4900 3100 -1900
rect 2300 -5000 3100 -4900
rect 9300 -1900 10100 -1800
rect 9300 -4900 9400 -1900
rect 10000 -4900 10100 -1900
rect 9300 -5000 10100 -4900
rect 14200 -1900 15000 -1800
rect 14200 -4900 14300 -1900
rect 14900 -4900 15000 -1900
rect 14200 -5000 15000 -4900
rect 20500 -1900 21300 -1800
rect 20500 -4900 20600 -1900
rect 21200 -4900 21300 -1900
rect 20500 -5000 21300 -4900
<< nsubdiff >>
rect -6900 3500 -6100 3600
rect -6900 500 -6800 3500
rect -6200 500 -6100 3500
rect -6900 400 -6100 500
rect -1500 3500 -700 3600
rect -1500 500 -1400 3500
rect -800 500 -700 3500
rect -1500 400 -700 500
rect 2400 3500 3200 3600
rect 2400 500 2500 3500
rect 3100 500 3200 3500
rect 2400 400 3200 500
rect 9200 3500 10000 3600
rect 9200 500 9300 3500
rect 9900 500 10000 3500
rect 9200 400 10000 500
rect 13100 3500 13900 3600
rect 13100 500 13200 3500
rect 13800 500 13900 3500
rect 13100 400 13900 500
rect 18500 3500 19300 3600
rect 18500 500 18600 3500
rect 19200 500 19300 3500
rect 18500 400 19300 500
<< psubdiffcont >>
rect -8800 -4900 -8200 -1900
rect -2500 -4900 -1900 -1900
rect 2400 -4900 3000 -1900
rect 9400 -4900 10000 -1900
rect 14300 -4900 14900 -1900
rect 20600 -4900 21200 -1900
<< nsubdiffcont >>
rect -6800 500 -6200 3500
rect -1400 500 -800 3500
rect 2500 500 3100 3500
rect 9300 500 9900 3500
rect 13200 500 13800 3500
rect 18600 500 19200 3500
<< poly >>
rect -5200 4050 -4800 4100
rect -5200 3750 -5150 4050
rect -4850 3750 -4800 4050
rect -5200 3600 -4800 3750
rect -3800 3700 16200 4100
rect -3800 3600 -3400 3700
rect -3300 3600 -2900 3700
rect 200 3600 600 3700
rect 700 3600 1100 3700
rect 4100 3600 4500 3700
rect 4600 3600 5000 3700
rect 7400 3600 7800 3700
rect 7900 3600 8300 3700
rect 11300 3600 11700 3700
rect 11800 3600 12200 3700
rect 15300 3600 15700 3700
rect 15800 3600 16200 3700
rect 17200 4050 17600 4100
rect 17200 3750 17250 4050
rect 17550 3750 17600 4050
rect 17200 3600 17600 3750
rect -5200 300 -4800 400
rect -3800 300 -3400 400
rect -3300 300 -2900 400
rect 200 300 600 400
rect 700 300 1100 400
rect 4100 300 4500 400
rect 4600 300 5000 400
rect 7400 300 7800 400
rect 7900 300 8300 400
rect 11300 300 11700 400
rect 11800 300 12200 400
rect 15300 300 15700 400
rect 15800 300 16200 400
rect 17200 300 17600 400
rect -5800 -1250 -3500 -1200
rect -7200 -1350 -6800 -1300
rect -7200 -1650 -7150 -1350
rect -6850 -1650 -6800 -1350
rect -7200 -1800 -6800 -1650
rect -5800 -1550 -3850 -1250
rect -3550 -1550 -3500 -1250
rect -5800 -1600 -3500 -1550
rect -900 -1250 4400 -1200
rect -900 -1550 1250 -1250
rect 1550 -1550 4400 -1250
rect -900 -1600 4400 -1550
rect -5800 -1800 -5400 -1600
rect -4400 -1800 -4000 -1700
rect -900 -1800 -500 -1600
rect 500 -1800 900 -1700
rect 4000 -1800 4400 -1600
rect 8000 -1250 13300 -1200
rect 8000 -1550 10850 -1250
rect 11150 -1550 13300 -1250
rect 8000 -1600 13300 -1550
rect 15900 -1250 18200 -1200
rect 15900 -1550 15950 -1250
rect 16250 -1550 18200 -1250
rect 15900 -1600 18200 -1550
rect 4500 -1800 4900 -1700
rect 7500 -1800 7900 -1700
rect 8000 -1800 8400 -1600
rect 11500 -1800 11900 -1700
rect 12900 -1800 13300 -1600
rect 16400 -1800 16800 -1700
rect 17800 -1800 18200 -1600
rect 19200 -1350 19600 -1300
rect 19200 -1650 19250 -1350
rect 19550 -1650 19600 -1350
rect 19200 -1800 19600 -1650
rect -7200 -5100 -6800 -5000
rect -5800 -5100 -5400 -5000
rect -4400 -5350 -4000 -5000
rect -900 -5100 -500 -5000
rect -4400 -5650 -4350 -5350
rect -4050 -5650 -4000 -5350
rect -4400 -5700 -4000 -5650
rect 500 -5350 900 -5000
rect 4000 -5100 4400 -5000
rect 500 -5650 550 -5350
rect 850 -5650 900 -5350
rect 500 -5700 900 -5650
rect 4500 -5350 4900 -5000
rect 7500 -5100 7900 -5000
rect 4500 -5650 4550 -5350
rect 4850 -5650 4900 -5350
rect 4500 -5700 4900 -5650
rect 8000 -5350 8400 -5000
rect 8000 -5650 8050 -5350
rect 8350 -5650 8400 -5350
rect 8000 -5700 8400 -5650
rect 11500 -5350 11900 -5000
rect 12900 -5100 13300 -5000
rect 11500 -5650 11550 -5350
rect 11850 -5650 11900 -5350
rect 11500 -5700 11900 -5650
rect 16400 -5350 16800 -5000
rect 17800 -5100 18200 -5000
rect 19200 -5100 19600 -5000
rect 16400 -5650 16450 -5350
rect 16750 -5650 16800 -5350
rect 16400 -5700 16800 -5650
<< polycont >>
rect -5150 3750 -4850 4050
rect 17250 3750 17550 4050
rect -7150 -1650 -6850 -1350
rect -3850 -1550 -3550 -1250
rect 1250 -1550 1550 -1250
rect 10850 -1550 11150 -1250
rect 15950 -1550 16250 -1250
rect 19250 -1650 19550 -1350
rect -4350 -5650 -4050 -5350
rect 550 -5650 850 -5350
rect 4550 -5650 4850 -5350
rect 8050 -5650 8350 -5350
rect 11550 -5650 11850 -5350
rect 16450 -5650 16750 -5350
<< locali >>
rect -5700 4050 -4800 4100
rect -5700 3750 -5150 4050
rect -4850 3750 -4800 4050
rect -5700 3700 -4800 3750
rect -5700 3600 -5300 3700
rect 6000 3600 6400 4800
rect 17200 4050 18100 4100
rect 17200 3750 17250 4050
rect 17550 3750 18100 4050
rect 17200 3700 18100 3750
rect 17700 3600 18100 3700
rect -6900 3500 -5300 3600
rect -6900 500 -6800 3500
rect -6200 500 -6000 3500
rect -5400 500 -5300 3500
rect -6900 400 -5300 500
rect -4700 3500 -3900 3600
rect -4700 500 -4600 3500
rect -4000 500 -3900 3500
rect -4700 400 -3900 500
rect -2800 3500 -2000 3600
rect -2800 500 -2700 3500
rect -2100 500 -2000 3500
rect -2800 400 -2000 500
rect -1500 3500 100 3600
rect -1500 500 -1400 3500
rect -800 500 -600 3500
rect 0 500 100 3500
rect -1500 400 100 500
rect 1200 3500 2000 3600
rect 1200 500 1300 3500
rect 1900 500 2000 3500
rect 1200 400 2000 500
rect 2400 3500 4000 3600
rect 2400 500 2500 3500
rect 3100 500 3300 3500
rect 3900 500 4000 3500
rect 2400 400 4000 500
rect 5100 3500 7300 3600
rect 5100 500 5200 3500
rect 5800 3200 6600 3500
rect 5800 500 5900 3200
rect 5100 400 5900 500
rect -5100 -650 -4700 -600
rect -5100 -950 -5050 -650
rect -4750 -950 -4700 -650
rect -7700 -1350 -6800 -1300
rect -7700 -1650 -7150 -1350
rect -6850 -1650 -6800 -1350
rect -7700 -1700 -6800 -1650
rect -7700 -1800 -7300 -1700
rect -5100 -1800 -4700 -950
rect -2800 -1000 -2400 400
rect -200 50 200 100
rect -200 -250 -150 50
rect 150 -250 200 50
rect -3900 -1250 -2400 -1200
rect -3900 -1550 -3850 -1250
rect -3550 -1550 -2400 -1250
rect -3900 -1600 -2400 -1550
rect -3900 -1800 -3500 -1600
rect -200 -1800 200 -250
rect 1200 -1000 1600 400
rect 1200 -1250 1600 -1200
rect 1200 -1550 1250 -1250
rect 1550 -1550 1600 -1250
rect 1200 -1800 1600 -1550
rect 6000 -1800 6400 3200
rect 6500 500 6600 3200
rect 7200 500 7300 3500
rect 6500 400 7300 500
rect 8400 3500 10000 3600
rect 8400 500 8500 3500
rect 9100 500 9300 3500
rect 9900 500 10000 3500
rect 8400 400 10000 500
rect 10400 3500 11200 3600
rect 10400 500 10500 3500
rect 11100 500 11200 3500
rect 10400 400 11200 500
rect 12300 3500 13900 3600
rect 12300 500 12400 3500
rect 13000 500 13200 3500
rect 13800 500 13900 3500
rect 12300 400 13900 500
rect 14400 3500 15200 3600
rect 14400 500 14500 3500
rect 15100 500 15200 3500
rect 14400 400 15200 500
rect 16300 3500 17100 3600
rect 16300 500 16400 3500
rect 17000 500 17100 3500
rect 16300 400 17100 500
rect 17700 3500 19300 3600
rect 17700 500 17800 3500
rect 18400 500 18600 3500
rect 19200 500 19300 3500
rect 17700 400 19300 500
rect 10800 -1250 11200 400
rect 10800 -1550 10850 -1250
rect 11150 -1550 11200 -1250
rect 10800 -1800 11200 -1550
rect 12200 50 12600 100
rect 12200 -250 12250 50
rect 12550 -250 12600 50
rect 12200 -1800 12600 -250
rect 14800 -1200 15200 400
rect 17100 -650 17500 -600
rect 17100 -950 17150 -650
rect 17450 -950 17500 -650
rect 14800 -1250 16300 -1200
rect 14800 -1550 15950 -1250
rect 16250 -1550 16300 -1250
rect 14800 -1600 16300 -1550
rect 15900 -1800 16300 -1600
rect 17100 -1800 17500 -950
rect 19200 -1350 20100 -1300
rect 19200 -1650 19250 -1350
rect 19550 -1650 20100 -1350
rect 19200 -1700 20100 -1650
rect 19700 -1800 20100 -1700
rect -8900 -1900 -7300 -1800
rect -8900 -4900 -8800 -1900
rect -8200 -4900 -8000 -1900
rect -7400 -4900 -7300 -1900
rect -8900 -5000 -7300 -4900
rect -6700 -1900 -5900 -1800
rect -6700 -4900 -6600 -1900
rect -6000 -4900 -5900 -1900
rect -6700 -5000 -5900 -4900
rect -5300 -1900 -4500 -1800
rect -5300 -4900 -5200 -1900
rect -4600 -4900 -4500 -1900
rect -5300 -5000 -4500 -4900
rect -3900 -1900 -3100 -1800
rect -3900 -4900 -3800 -1900
rect -3200 -4900 -3100 -1900
rect -3900 -5000 -3100 -4900
rect -2600 -1900 -1000 -1800
rect -2600 -4900 -2500 -1900
rect -1900 -4900 -1700 -1900
rect -1100 -4900 -1000 -1900
rect -2600 -5000 -1000 -4900
rect -400 -1900 400 -1800
rect -400 -4900 -300 -1900
rect 300 -4900 400 -1900
rect -400 -5000 400 -4900
rect 1000 -1900 1800 -1800
rect 1000 -4900 1100 -1900
rect 1700 -4900 1800 -1900
rect 1000 -5000 1800 -4900
rect 2300 -1900 3900 -1800
rect 2300 -4900 2400 -1900
rect 3000 -4900 3200 -1900
rect 3800 -4900 3900 -1900
rect 2300 -5000 3900 -4900
rect 5000 -1900 7400 -1800
rect 5000 -4900 5100 -1900
rect 5700 -2200 6700 -1900
rect 5700 -4900 5800 -2200
rect 5000 -5000 5800 -4900
rect 6600 -4900 6700 -2200
rect 7300 -4900 7400 -1900
rect 6600 -5000 7400 -4900
rect 8500 -1900 10100 -1800
rect 8500 -4900 8600 -1900
rect 9200 -4900 9400 -1900
rect 10000 -4900 10100 -1900
rect 8500 -5000 10100 -4900
rect 10600 -1900 11400 -1800
rect 10600 -4900 10700 -1900
rect 11300 -4900 11400 -1900
rect 10600 -5000 11400 -4900
rect 12000 -1900 12800 -1800
rect 12000 -4900 12100 -1900
rect 12700 -4900 12800 -1900
rect 12000 -5000 12800 -4900
rect 13400 -1900 15000 -1800
rect 13400 -4900 13500 -1900
rect 14100 -4900 14300 -1900
rect 14900 -4900 15000 -1900
rect 13400 -5000 15000 -4900
rect 15500 -1900 16300 -1800
rect 15500 -4900 15600 -1900
rect 16200 -4900 16300 -1900
rect 15500 -5000 16300 -4900
rect 16900 -1900 17700 -1800
rect 16900 -4900 17000 -1900
rect 17600 -4900 17700 -1900
rect 16900 -5000 17700 -4900
rect 18300 -1900 19100 -1800
rect 18300 -4900 18400 -1900
rect 19000 -4900 19100 -1900
rect 18300 -5000 19100 -4900
rect 19700 -1900 21300 -1800
rect 19700 -4900 19800 -1900
rect 20400 -4900 20600 -1900
rect 21200 -4900 21300 -1900
rect 19700 -5000 21300 -4900
rect -4400 -5350 -4000 -5300
rect -4400 -5650 -4350 -5350
rect -4050 -5650 -4000 -5350
rect -4400 -5700 -4000 -5650
rect 500 -5350 900 -5300
rect 500 -5650 550 -5350
rect 850 -5650 900 -5350
rect 500 -5700 900 -5650
rect 4500 -5350 4900 -5300
rect 4500 -5650 4550 -5350
rect 4850 -5650 4900 -5350
rect 4500 -5700 4900 -5650
rect 8000 -5350 8400 -5300
rect 8000 -5650 8050 -5350
rect 8350 -5650 8400 -5350
rect 8000 -5700 8400 -5650
rect 11500 -5350 11900 -5300
rect 11500 -5650 11550 -5350
rect 11850 -5650 11900 -5350
rect 11500 -5700 11900 -5650
rect 16400 -5350 16800 -5300
rect 16400 -5650 16450 -5350
rect 16750 -5650 16800 -5350
rect 16400 -5700 16800 -5650
<< viali >>
rect -6800 500 -6200 3500
rect -6000 500 -5400 3500
rect -4600 500 -4000 3500
rect -1400 500 -800 3500
rect -600 500 0 3500
rect 2500 500 3100 3500
rect 3300 500 3900 3500
rect -5050 -950 -4750 -650
rect -150 -250 150 50
rect 8500 500 9100 3500
rect 9300 500 9900 3500
rect 12400 500 13000 3500
rect 13200 500 13800 3500
rect 16400 500 17000 3500
rect 17800 500 18400 3500
rect 18600 500 19200 3500
rect 12250 -250 12550 50
rect 17150 -950 17450 -650
rect -8800 -4900 -8200 -1900
rect -8000 -4900 -7400 -1900
rect -6600 -4900 -6000 -1900
rect -2500 -4900 -1900 -1900
rect -1700 -4900 -1100 -1900
rect 2400 -4900 3000 -1900
rect 3200 -4900 3800 -1900
rect 8600 -4900 9200 -1900
rect 9400 -4900 10000 -1900
rect 13500 -4900 14100 -1900
rect 14300 -4900 14900 -1900
rect 18400 -4900 19000 -1900
rect 19800 -4900 20400 -1900
rect 20600 -4900 21200 -1900
rect -4350 -5650 -4050 -5350
rect 550 -5650 850 -5350
rect 4550 -5650 4850 -5350
rect 8050 -5650 8350 -5350
rect 11550 -5650 11850 -5350
rect 16450 -5650 16750 -5350
<< metal1 >>
rect -8900 3500 19300 3600
rect -8900 500 -6800 3500
rect -6200 500 -6000 3500
rect -5400 500 -4600 3500
rect -4000 500 -1400 3500
rect -800 500 -600 3500
rect 0 500 2500 3500
rect 3100 500 3300 3500
rect 3900 500 8500 3500
rect 9100 500 9300 3500
rect 9900 500 12400 3500
rect 13000 500 13200 3500
rect 13800 500 16400 3500
rect 17000 500 17800 3500
rect 18400 500 18600 3500
rect 19200 500 19300 3500
rect -8900 400 19300 500
rect -8900 50 12600 100
rect -8900 -250 -150 50
rect 150 -250 12250 50
rect 12550 -250 12600 50
rect -8900 -300 12600 -250
rect -8900 -650 17500 -600
rect -8900 -950 -5050 -650
rect -4750 -950 17150 -650
rect 17450 -950 17500 -650
rect -8900 -1000 17500 -950
rect -8900 -1900 21300 -1800
rect -8900 -4900 -8800 -1900
rect -8200 -4900 -8000 -1900
rect -7400 -4900 -6600 -1900
rect -6000 -4900 -2500 -1900
rect -1900 -4900 -1700 -1900
rect -1100 -4900 2400 -1900
rect 3000 -4900 3200 -1900
rect 3800 -4900 8600 -1900
rect 9200 -4900 9400 -1900
rect 10000 -4900 13500 -1900
rect 14100 -4900 14300 -1900
rect 14900 -4900 18400 -1900
rect 19000 -4900 19800 -1900
rect 20400 -4900 20600 -1900
rect 21200 -4900 21300 -1900
rect -8900 -5000 21300 -4900
rect -8900 -5350 16800 -5300
rect -8900 -5650 -4350 -5350
rect -4050 -5650 550 -5350
rect 850 -5650 4550 -5350
rect 4850 -5650 8050 -5350
rect 8350 -5650 11550 -5350
rect 11850 -5650 16450 -5350
rect 16750 -5650 16800 -5350
rect -8900 -5700 16800 -5650
<< labels >>
flabel locali 6200 4800 6200 4800 0 FreeSans 4000 0 0 0 i_fvf_out
flabel metal1 -8900 2100 -8900 2100 0 FreeSans 4000 0 0 0 VP
flabel metal1 -8900 -100 -8900 -100 0 FreeSans 4000 0 0 0 i_out
flabel metal1 -8900 -800 -8900 -800 0 FreeSans 4000 0 0 0 i_dump
flabel metal1 -8900 -3400 -8900 -3400 0 FreeSans 4000 0 0 0 VN
flabel metal1 -8900 -5500 -8900 -5500 0 FreeSans 4000 0 0 0 VCN
<< end >>
