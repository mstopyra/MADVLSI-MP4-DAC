magic
tech sky130A
magscale 1 2
timestamp 1701235168
<< error_p >>
rect -60000 -20800 -59800 -15860
rect -59000 -20800 -58983 -15860
rect -51817 -20800 -51800 -15860
rect -44017 -20800 -44000 -15860
rect -43200 -20800 -41400 -15860
<< poly >>
rect 9400 -11700 10200 -11600
rect 9400 -12200 9500 -11700
rect 7200 -12300 9500 -12200
rect 10100 -12300 10200 -11700
rect 7200 -12400 10200 -12300
<< polycont >>
rect 9500 -12300 10100 -11700
<< locali >>
rect 9400 -11700 10200 -11600
rect 9400 -12300 9500 -11700
rect 10100 -12300 10200 -11700
rect 9400 -12400 10200 -12300
rect -7100 -19800 -5900 -19600
rect -7100 -32200 -6300 -19800
rect -20400 -33000 -6300 -32200
<< viali >>
rect -34900 37900 -34700 38100
rect 9500 -12300 10100 -11700
rect -41100 -24700 -40500 -24100
<< metal1 >>
rect -35000 38100 -34600 38200
rect -35000 37900 -34900 38100
rect -34700 37900 -34600 38100
rect -35000 37800 -34600 37900
rect -58000 28000 -57200 28100
rect -58000 27400 -57900 28000
rect -57300 27400 -57200 28000
rect -58000 24200 -57200 27400
rect -60200 17800 -52400 24200
rect -58000 17000 -52700 17800
rect -42000 16800 -34000 23200
rect -2400 15800 17800 22200
rect -96000 0 -59800 2400
rect -58000 0 -36400 2200
rect -32000 0 -4000 2200
rect -96000 -10000 9200 0
rect -96000 -12200 -74400 -10000
rect -71000 -14600 -14600 -10000
rect -6000 -12600 9200 -10000
rect 9400 -11700 10200 -11600
rect 9400 -12300 9500 -11700
rect 10100 -12300 10200 -11700
rect 9400 -12400 10200 -12300
rect 11400 -20400 17800 15800
rect -41200 -24100 -40400 -24000
rect -41200 -24700 -41100 -24100
rect -40500 -24700 -40400 -24100
rect -41200 -24800 -40400 -24700
rect -10600 -31600 -6000 -20400
rect 9000 -26800 17800 -20400
rect 11400 -34700 17800 -26800
rect -80000 -41100 17800 -34700
<< via1 >>
rect -34900 37900 -34700 38100
rect -57900 27400 -57300 28000
rect 9500 -12300 10100 -11700
rect -33700 -22100 -33100 -21500
rect -18900 -23500 -18300 -22900
rect -41100 -24700 -40500 -24100
<< metal2 >>
rect -36400 38100 -34600 38200
rect -36400 37900 -34900 38100
rect -34700 37900 -34600 38100
rect -36400 37800 -34600 37900
rect -36400 27300 -35700 37800
rect 2800 32000 4400 32800
rect -58000 17000 -57200 24600
rect -77000 16400 -57200 17000
rect -79600 1700 -78800 1900
rect -79600 1100 -79500 1700
rect -78900 1100 -78800 1700
rect -79600 1000 -78800 1100
rect -33800 -21500 -33000 27200
rect -33800 -22100 -33700 -21500
rect -33100 -22100 -33000 -21500
rect -33800 -22200 -33000 -22100
rect 3600 -22800 4400 32000
rect -19000 -22900 4400 -22800
rect -19000 -23500 -18900 -22900
rect -18300 -23500 4400 -22900
rect -19000 -23600 4400 -23500
rect 9400 -11700 10200 -11600
rect 9400 -12300 9500 -11700
rect 10100 -12300 10200 -11700
rect -74300 -24100 -40400 -24000
rect -74300 -24700 -41100 -24100
rect -40500 -24700 -40400 -24100
rect -74300 -24800 -40400 -24700
rect -74300 -30600 -73500 -24800
rect 9400 -33300 10200 -12300
rect -75100 -34100 10200 -33300
<< via2 >>
rect -79500 1100 -78900 1700
<< metal3 >>
rect -79600 1700 -72700 1800
rect -79600 1100 -79500 1700
rect -78900 1100 -72700 1700
rect -79600 1000 -72700 1100
rect -73500 -34100 -72700 1000
use 7BIT_DAC_block  7BIT_DAC_block_0
timestamp 1701150204
transform 1 0 -39000 0 1 2200
box 4000 -200 41800 36000
use BIASGEN_VBP_VBN  BIASGEN_VBP_VBN_0
timestamp 1701228322
transform 1 0 -94600 0 -1 24201
box -1400 -600 34800 22400
use first_current_mirror  first_current_mirror_0
timestamp 1701232898
transform 1 0 -55500 0 1 2900
box -2500 -900 19100 43100
use FVF_block  FVF_block_0
timestamp 1701232898
transform 1 0 -53200 0 1 -21600
box -17800 -11400 42800 9600
use REAL_VCN_BIAS_GEN  REAL_VCN_BIAS_GEN_0
timestamp 1701222951
transform 1 0 -3200 0 1 -33200
box -2800 5800 12400 21200
use second_current_mirror  second_current_mirror_0
timestamp 1701228322
transform -1 0 -76774 0 1 -55000
box -2500 -800 19100 43000
<< end >>
