magic
tech sky130A
timestamp 1701117479
<< nwell >>
rect -400 800 1100 7400
<< nmos >>
rect 300 7700 700 10900
<< pmos >>
rect 300 900 700 7300
<< ndiff >>
rect 0 10800 300 10900
rect 0 7800 100 10800
rect 200 7800 300 10800
rect 0 7700 300 7800
rect 700 10800 1000 10900
rect 700 7800 800 10800
rect 900 7800 1000 10800
rect 700 7700 1000 7800
<< pdiff >>
rect 0 7200 300 7300
rect 0 1000 100 7200
rect 200 1000 300 7200
rect 0 900 300 1000
rect 700 7200 1000 7300
rect 700 1000 800 7200
rect 900 1000 1000 7200
rect 700 900 1000 1000
<< ndiffc >>
rect 100 7800 200 10800
rect 800 7800 900 10800
<< pdiffc >>
rect 100 1000 200 7200
rect 800 1000 900 7200
<< psubdiff >>
rect -300 10800 0 10900
rect -300 7800 -200 10800
rect -100 7800 0 10800
rect -300 7700 0 7800
<< nsubdiff >>
rect -300 7200 0 7300
rect -300 1000 -200 7200
rect -100 1000 0 7200
rect -300 900 0 1000
<< psubdiffcont >>
rect -200 7800 -100 10800
<< nsubdiffcont >>
rect -200 1000 -100 7200
<< poly >>
rect 300 10900 700 11000
rect 300 7550 700 7700
rect 300 7450 350 7550
rect 650 7450 700 7550
rect 300 7300 700 7450
rect 300 800 700 900
<< polycont >>
rect 350 7450 650 7550
<< locali >>
rect -300 10800 200 10900
rect -300 7800 -200 10800
rect -100 7800 100 10800
rect -300 7700 200 7800
rect 700 10800 1000 10900
rect 700 7800 800 10800
rect 900 7800 1000 10800
rect 700 7700 1000 7800
rect 300 7550 700 7600
rect 900 7550 1000 7700
rect 200 7450 350 7550
rect 650 7450 800 7550
rect 900 7450 1100 7550
rect 300 7400 700 7450
rect 900 7300 1000 7450
rect -300 7200 200 7300
rect -300 1000 -200 7200
rect -100 1000 100 7200
rect -300 900 200 1000
rect 700 7200 1000 7300
rect 700 1000 800 7200
rect 900 1000 1000 7200
rect 700 900 1000 1000
<< viali >>
rect -200 7800 -100 10800
rect 100 7800 200 10800
rect -200 1000 -100 7200
rect 100 1000 200 7200
<< metal1 >>
rect -400 10800 1000 10900
rect -400 7800 -200 10800
rect -100 7800 100 10800
rect 200 7800 1000 10800
rect -400 7700 1000 7800
rect -400 7200 1000 7300
rect -400 1000 -200 7200
rect -100 1000 100 7200
rect 200 1000 1000 7200
rect -400 900 1000 1000
<< labels >>
flabel metal1 -400 5700 -400 5700 7 FreeSans 800 0 0 0 VP
port 3 w
flabel metal1 -400 9700 -400 9700 7 FreeSans 800 0 0 0 VN
port 4 w
flabel locali 1100 7500 1100 7500 3 FreeSans 800 0 0 0 Q
port 6 e
flabel poly 500 800 500 800 5 FreeSans 800 0 0 0 A
port 5 s
<< end >>
