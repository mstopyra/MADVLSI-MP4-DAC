* NGSPICE file created from 7BIT_DAC_block.ext - technology: sky130A

X0 DAC_block_20/inverter_0/Q DAC_block_20/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X1 DAC_block_20/inverter_0/Q DAC_block_20/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=192 ps=134 w=64 l=4
X2 I_DUMP DAC_block_20/inverter_0/Q DAC_block_20/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X3 DAC_block_20/a_5400_7600# I_IN DAC_block_20/H_V VN sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X4 DAC_block_15/H_V I_IN DAC_block_20/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X5 DAC_block_20/H_V DAC_block_20/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X6 DAC_block_14/inverter_0/Q DAC_block_14/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=939 ps=686 w=32 l=4
X7 DAC_block_14/inverter_0/Q DAC_block_14/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=903 ps=644 w=64 l=4
X8 I_DUMP DAC_block_14/inverter_0/Q DAC_block_14/H_V VN sky130_fd_pr__nfet_01v8 ad=768 pd=560 as=279 ps=201 w=32 l=4
X9 DAC_block_14/a_5400_7600# I_IN DAC_block_14/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X10 DAC_block_16/H_V I_IN DAC_block_14/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=288 pd=210 as=0 ps=0 w=32 l=4
X11 DAC_block_14/H_V DAC_block_14/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=837 ps=609 w=32 l=4
X12 DAC_block_15/inverter_0/Q DAC_block_15/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=0 ps=0 w=32 l=4
X13 DAC_block_15/inverter_0/Q DAC_block_15/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=0 ps=0 w=64 l=4
X14 I_DUMP DAC_block_15/inverter_0/Q DAC_block_15/H_V VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=288 ps=210 w=32 l=4
X15 DAC_block_15/a_5400_7600# I_IN DAC_block_15/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X16 DAC_block_15/H_V_OUT I_IN DAC_block_15/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=258 pd=177 as=0 ps=0 w=32 l=4
X17 DAC_block_15/H_V DAC_block_15/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X18 DAC_block_16/inverter_0/Q DAC_block_16/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=0 ps=0 w=32 l=4
X19 DAC_block_16/inverter_0/Q DAC_block_16/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=0 ps=0 w=64 l=4
X20 I_DUMP DAC_block_16/inverter_0/Q DAC_block_16/H_V VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X21 DAC_block_16/a_5400_7600# I_IN DAC_block_16/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X22 DAC_block_17/H_V I_IN DAC_block_16/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=288 pd=210 as=0 ps=0 w=32 l=4
X23 DAC_block_16/H_V DAC_block_16/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X24 DAC_block_17/inverter_0/Q DAC_block_17/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=0 ps=0 w=32 l=4
X25 DAC_block_17/inverter_0/Q DAC_block_17/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=0 ps=0 w=64 l=4
X26 I_DUMP DAC_block_17/inverter_0/Q DAC_block_17/H_V VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X27 DAC_block_17/a_5400_7600# I_IN DAC_block_17/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X28 DAC_block_18/H_V I_IN DAC_block_17/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=288 pd=210 as=0 ps=0 w=32 l=4
X29 DAC_block_17/H_V DAC_block_17/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X30 DAC_block_18/inverter_0/Q DAC_block_18/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=0 ps=0 w=32 l=4
X31 DAC_block_18/inverter_0/Q DAC_block_18/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=0 ps=0 w=64 l=4
X32 I_DUMP DAC_block_18/inverter_0/Q DAC_block_18/H_V VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X33 DAC_block_18/a_5400_7600# I_IN DAC_block_18/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X34 DAC_block_19/H_V I_IN DAC_block_18/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=288 pd=210 as=0 ps=0 w=32 l=4
X35 DAC_block_18/H_V DAC_block_18/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X36 DAC_block_19/inverter_0/Q DAC_block_19/D_IN VN VN sky130_fd_pr__nfet_01v8 ad=105 pd=79 as=0 ps=0 w=32 l=4
X37 DAC_block_19/inverter_0/Q DAC_block_19/D_IN DAC_block_20/VP DAC_block_20/VP sky130_fd_pr__pfet_01v8 ad=192 pd=134 as=0 ps=0 w=64 l=4
X38 I_DUMP DAC_block_19/inverter_0/Q DAC_block_19/H_V VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X39 DAC_block_19/a_5400_7600# I_IN DAC_block_19/H_V VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=0 ps=0 w=32 l=4
X40 DAC_block_20/H_V I_IN DAC_block_19/a_5400_7600# VN sky130_fd_pr__nfet_01v8 ad=288 pd=210 as=0 ps=0 w=32 l=4
X41 DAC_block_19/H_V DAC_block_19/D_IN I_OUT VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=32 l=4
X42 I_DUMP I_IN DAC_block_15/H_V_OUT VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X43 I_OUT VN VN VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X44 I_OUT VN VN VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X45 DAC_block_14/H_V VN VN VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X46 DAC_block_15/H_V_OUT VN VN VN sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
