magic
tech sky130A
timestamp 1701221553
<< nwell >>
rect -1400 7000 6100 10600
<< nmos >>
rect -1100 3200 -700 6400
rect -400 3200 0 6400
rect 100 3200 500 6400
rect 600 3200 1000 6400
rect 1100 3200 1500 6400
rect 1800 3200 2200 6400
rect 2500 3200 2900 6400
rect 3200 3200 3600 6400
rect 3700 3200 4100 6400
rect 4200 3200 4600 6400
rect 4700 3200 5100 6400
rect 5400 3200 5800 6400
<< pmos >>
rect -1100 7100 -700 10300
rect -400 7100 0 10300
rect 100 7100 500 10300
rect 600 7100 1000 10300
rect 1100 7100 1500 10300
rect 1600 7100 2000 10300
rect 2300 7100 2700 10300
rect 2800 7100 3200 10300
rect 3300 7100 3700 10300
rect 3800 7100 4200 10300
rect 4300 7100 4700 10300
rect 5000 7100 5400 10300
<< ndiff >>
rect -1200 6380 -1100 6400
rect -1200 3220 -1180 6380
rect -1120 3220 -1100 6380
rect -1200 3200 -1100 3220
rect -700 6380 -600 6400
rect -500 6380 -400 6400
rect -700 3220 -680 6380
rect -620 3220 -600 6380
rect -500 3220 -480 6380
rect -420 3220 -400 6380
rect -700 3200 -600 3220
rect -500 3200 -400 3220
rect 0 6380 100 6400
rect 0 3220 20 6380
rect 80 3220 100 6380
rect 0 3200 100 3220
rect 500 6380 600 6400
rect 500 3220 520 6380
rect 580 3220 600 6380
rect 500 3200 600 3220
rect 1000 6380 1100 6400
rect 1000 3220 1020 6380
rect 1080 3220 1100 6380
rect 1000 3200 1100 3220
rect 1500 6380 1600 6400
rect 1700 6380 1800 6400
rect 1500 3220 1520 6380
rect 1580 3220 1600 6380
rect 1700 3220 1720 6380
rect 1780 3220 1800 6380
rect 1500 3200 1600 3220
rect 1700 3200 1800 3220
rect 2200 6380 2500 6400
rect 2200 3220 2220 6380
rect 2480 3220 2500 6380
rect 2200 3200 2500 3220
rect 2900 6380 3000 6400
rect 3100 6380 3200 6400
rect 2900 3220 2920 6380
rect 2980 3220 3000 6380
rect 3100 3220 3120 6380
rect 3180 3220 3200 6380
rect 2900 3200 3000 3220
rect 3100 3200 3200 3220
rect 3600 6380 3700 6400
rect 3600 3220 3620 6380
rect 3680 3220 3700 6380
rect 3600 3200 3700 3220
rect 4100 6380 4200 6400
rect 4100 3220 4120 6380
rect 4180 3220 4200 6380
rect 4100 3200 4200 3220
rect 4600 6380 4700 6400
rect 4600 3220 4620 6380
rect 4680 3220 4700 6380
rect 4600 3200 4700 3220
rect 5100 6380 5200 6400
rect 5300 6380 5400 6400
rect 5100 3220 5120 6380
rect 5180 3220 5200 6380
rect 5300 3220 5320 6380
rect 5380 3220 5400 6380
rect 5100 3200 5200 3220
rect 5300 3200 5400 3220
rect 5800 6380 5900 6400
rect 5800 3220 5820 6380
rect 5880 3220 5900 6380
rect 5800 3200 5900 3220
<< pdiff >>
rect -1200 10280 -1100 10300
rect -1200 7120 -1180 10280
rect -1120 7120 -1100 10280
rect -1200 7100 -1100 7120
rect -700 10280 -600 10300
rect -500 10280 -400 10300
rect -700 7120 -680 10280
rect -620 7120 -600 10280
rect -500 7120 -480 10280
rect -420 7120 -400 10280
rect -700 7100 -600 7120
rect -500 7100 -400 7120
rect 0 7100 100 10300
rect 500 7100 600 10300
rect 1000 7100 1100 10300
rect 1500 7100 1600 10300
rect 2000 10280 2100 10300
rect 2200 10280 2300 10300
rect 2000 7120 2020 10280
rect 2080 7120 2100 10280
rect 2200 7120 2220 10280
rect 2280 7120 2300 10280
rect 2000 7100 2100 7120
rect 2200 7100 2300 7120
rect 2700 7100 2800 10300
rect 3200 7100 3300 10300
rect 3700 7100 3800 10300
rect 4200 7100 4300 10300
rect 4700 10280 4800 10300
rect 4900 10280 5000 10300
rect 4700 7120 4720 10280
rect 4780 7120 4800 10280
rect 4900 7120 4920 10280
rect 4980 7120 5000 10280
rect 4700 7100 4800 7120
rect 4900 7100 5000 7120
rect 5400 10280 5500 10300
rect 5400 7120 5420 10280
rect 5480 7120 5500 10280
rect 5400 7100 5500 7120
<< ndiffc >>
rect -1180 3220 -1120 6380
rect -680 3220 -620 6380
rect -480 3220 -420 6380
rect 20 3220 80 6380
rect 520 3220 580 6380
rect 1020 3220 1080 6380
rect 1520 3220 1580 6380
rect 1720 3220 1780 6380
rect 2220 3220 2480 6380
rect 2920 3220 2980 6380
rect 3120 3220 3180 6380
rect 3620 3220 3680 6380
rect 4120 3220 4180 6380
rect 4620 3220 4680 6380
rect 5120 3220 5180 6380
rect 5320 3220 5380 6380
rect 5820 3220 5880 6380
<< pdiffc >>
rect -1180 7120 -1120 10280
rect -680 7120 -620 10280
rect -480 7120 -420 10280
rect 2020 7120 2080 10280
rect 2220 7120 2280 10280
rect 4720 7120 4780 10280
rect 4920 7120 4980 10280
rect 5420 7120 5480 10280
<< psubdiff >>
rect -1300 6380 -1200 6400
rect -1300 3220 -1280 6380
rect -1220 3220 -1200 6380
rect -1300 3200 -1200 3220
rect -600 6380 -500 6400
rect -600 3220 -580 6380
rect -520 3220 -500 6380
rect -600 3200 -500 3220
rect 1600 6380 1700 6400
rect 1600 3220 1620 6380
rect 1680 3220 1700 6380
rect 1600 3200 1700 3220
rect 3000 6380 3100 6400
rect 3000 3220 3020 6380
rect 3080 3220 3100 6380
rect 3000 3200 3100 3220
rect 5200 6380 5300 6400
rect 5200 3220 5220 6380
rect 5280 3220 5300 6380
rect 5200 3200 5300 3220
rect 5900 6380 6000 6400
rect 5900 3220 5920 6380
rect 5980 3220 6000 6380
rect 5900 3200 6000 3220
<< nsubdiff >>
rect -600 10280 -500 10300
rect -600 7120 -580 10280
rect -520 7120 -500 10280
rect -600 7100 -500 7120
rect 2100 10280 2200 10300
rect 2100 7120 2120 10280
rect 2180 7120 2200 10280
rect 2100 7100 2200 7120
rect 4800 10280 4900 10300
rect 4800 7120 4820 10280
rect 4880 7120 4900 10280
rect 4800 7100 4900 7120
<< psubdiffcont >>
rect -1280 3220 -1220 6380
rect -580 3220 -520 6380
rect 1620 3220 1680 6380
rect 3020 3220 3080 6380
rect 5220 3220 5280 6380
rect 5920 3220 5980 6380
<< nsubdiffcont >>
rect -580 7120 -520 10280
rect 2120 7120 2180 10280
rect 4820 7120 4880 10280
<< poly >>
rect -1400 10400 5300 10500
rect -1000 10325 -800 10400
rect -300 10325 -100 10400
rect 200 10325 400 10400
rect 700 10325 900 10400
rect 1200 10325 1400 10400
rect 1700 10325 1900 10400
rect 2400 10325 2600 10400
rect 2900 10325 3100 10400
rect 3400 10325 3600 10400
rect 3900 10325 4100 10400
rect 4400 10325 4600 10400
rect 5100 10325 5300 10400
rect -1100 10300 -700 10325
rect -400 10300 0 10325
rect 100 10300 500 10325
rect 600 10300 1000 10325
rect 1100 10300 1500 10325
rect 1600 10300 2000 10325
rect 2300 10300 2700 10325
rect 2800 10300 3200 10325
rect 3300 10300 3700 10325
rect 3800 10300 4200 10325
rect 4300 10300 4700 10325
rect 5000 10300 5400 10325
rect -1100 7075 -700 7100
rect -400 7075 0 7100
rect 100 7075 500 7100
rect 600 7075 1000 7100
rect 1100 7075 1500 7100
rect 1600 7075 2000 7100
rect 2300 7075 2700 7100
rect 2800 7075 3200 7100
rect 3300 7075 3700 7100
rect 3800 7075 4200 7100
rect 4300 7075 4700 7100
rect 5000 7075 5400 7100
rect 2000 6980 2200 7000
rect 2000 6920 2120 6980
rect 2180 6920 2200 6980
rect 2000 6900 2200 6920
rect 2000 6700 2100 6900
rect -1200 6590 -1000 6600
rect -1200 6510 -1190 6590
rect -1110 6510 -1000 6590
rect -1200 6500 -1000 6510
rect -1100 6420 -1000 6500
rect 1200 6500 3500 6700
rect 1200 6420 1400 6500
rect 1900 6420 2100 6500
rect 2600 6420 2800 6500
rect 3300 6420 3500 6500
rect 5700 6590 5900 6600
rect 5700 6510 5810 6590
rect 5890 6510 5900 6590
rect 5700 6500 5900 6510
rect 5700 6420 5800 6500
rect -1100 6400 -700 6420
rect -400 6400 0 6420
rect 100 6400 500 6420
rect 600 6400 1000 6420
rect 1100 6400 1500 6420
rect 1800 6400 2200 6420
rect 2500 6400 2900 6420
rect 3200 6400 3600 6420
rect 3700 6400 4100 6420
rect 4200 6400 4600 6420
rect 4700 6400 5100 6420
rect 5400 6400 5800 6420
rect -1100 3180 -700 3200
rect -400 3180 0 3200
rect 100 3180 500 3200
rect 600 3180 1000 3200
rect 1100 3180 1500 3200
rect 1800 3180 2200 3200
rect 2500 3180 2900 3200
rect 3200 3180 3600 3200
rect 3700 3180 4100 3200
rect 4200 3180 4600 3200
rect 4700 3180 5100 3200
rect 5400 3180 5800 3200
rect -200 3050 0 3180
rect -200 2950 -150 3050
rect -50 2950 0 3050
rect -200 2900 0 2950
rect 200 3050 400 3180
rect 200 2950 250 3050
rect 350 2950 400 3050
rect 200 2900 400 2950
rect 700 3050 900 3180
rect 700 2950 750 3050
rect 850 2950 900 3050
rect 700 2900 900 2950
rect 1100 3050 1300 3180
rect 1100 2950 1150 3050
rect 1250 2950 1300 3050
rect 1100 2900 1300 2950
rect 3400 3050 3600 3180
rect 3400 2950 3450 3050
rect 3550 2950 3600 3050
rect 3400 2900 3600 2950
rect 3800 3050 4000 3180
rect 3800 2950 3850 3050
rect 3950 2950 4000 3050
rect 3800 2900 4000 2950
rect 4300 3050 4500 3180
rect 4300 2950 4350 3050
rect 4450 2950 4500 3050
rect 4300 2900 4500 2950
rect 4700 3050 4900 3180
rect 4700 2950 4750 3050
rect 4850 2950 4900 3050
rect 4700 2900 4900 2950
<< polycont >>
rect 2120 6920 2180 6980
rect -1190 6510 -1110 6590
rect 5810 6510 5890 6590
rect -150 2950 -50 3050
rect 250 2950 350 3050
rect 750 2950 850 3050
rect 1150 2950 1250 3050
rect 3450 2950 3550 3050
rect 3850 2950 3950 3050
rect 4350 2950 4450 3050
rect 4750 2950 4850 3050
<< locali >>
rect -1190 10280 -1110 10300
rect -1190 7120 -1180 10280
rect -1120 7120 -1110 10280
rect -1190 7000 -1110 7120
rect -690 10280 -610 10300
rect -690 7120 -680 10280
rect -620 7120 -610 10280
rect -690 7100 -610 7120
rect -590 10280 -510 10300
rect -590 7120 -580 10280
rect -520 7120 -510 10280
rect -590 7100 -510 7120
rect -490 10280 -410 10300
rect -490 7120 -480 10280
rect -420 7120 -410 10280
rect -490 7110 -410 7120
rect 2010 10280 2090 10300
rect 2010 7120 2020 10280
rect 2080 7120 2090 10280
rect 2010 7080 2090 7120
rect 2110 10280 2190 10300
rect 2110 7120 2120 10280
rect 2180 7120 2190 10280
rect 2110 7100 2190 7120
rect 2210 10280 2290 10300
rect 2210 7120 2220 10280
rect 2280 7120 2290 10280
rect 2210 7080 2290 7120
rect 4710 10290 4790 10300
rect 4910 10290 4990 10300
rect 4710 10280 4990 10290
rect 4710 7120 4720 10280
rect 4780 7120 4820 10280
rect 4880 7120 4920 10280
rect 4980 7120 4990 10280
rect 4710 7110 4990 7120
rect 5410 10280 5490 10300
rect 5410 7120 5420 10280
rect 5480 7120 5490 10280
rect 2010 7000 2290 7080
rect 5410 7000 5490 7120
rect -1200 6800 -1100 7000
rect 2100 6980 2200 7000
rect 2100 6920 2120 6980
rect 2180 6920 2200 6980
rect 2100 6900 2200 6920
rect 5400 6800 5500 7000
rect -1400 6700 5900 6800
rect -1200 6590 -1100 6700
rect -1200 6510 -1190 6590
rect -1110 6510 -1100 6590
rect -1200 6500 -1100 6510
rect -700 6500 5400 6600
rect 5800 6590 5900 6700
rect 5800 6510 5810 6590
rect 5890 6510 5900 6590
rect 5800 6500 5900 6510
rect -1290 6380 -1210 6390
rect -1290 3220 -1280 6380
rect -1220 3220 -1210 6380
rect -1290 3210 -1210 3220
rect -1190 6380 -1110 6500
rect -1190 3220 -1180 6380
rect -1120 3220 -1110 6380
rect -1190 3210 -1110 3220
rect -690 6380 -610 6500
rect -690 3220 -680 6380
rect -620 3220 -610 6380
rect -690 3210 -610 3220
rect -590 6380 -510 6390
rect -590 3220 -580 6380
rect -520 3220 -510 6380
rect -590 3210 -510 3220
rect -490 6380 -410 6500
rect -490 3220 -480 6380
rect -420 3220 -410 6380
rect -490 3200 -410 3220
rect 10 6380 90 6390
rect 10 3220 20 6380
rect 80 3220 90 6380
rect 10 3100 90 3220
rect 510 6380 590 6390
rect 510 3220 520 6380
rect 580 3220 590 6380
rect 510 3100 590 3220
rect 1010 6380 1090 6390
rect 1010 3220 1020 6380
rect 1080 3220 1090 6380
rect 1010 3100 1090 3220
rect 1510 6380 1590 6500
rect 1510 3220 1520 6380
rect 1580 3220 1590 6380
rect 1510 3200 1590 3220
rect 1610 6380 1690 6390
rect 1610 3220 1620 6380
rect 1680 3220 1690 6380
rect 1610 3210 1690 3220
rect 1710 6380 1790 6500
rect 1710 3220 1720 6380
rect 1780 3220 1790 6380
rect 1710 3210 1790 3220
rect 2200 6380 2500 6400
rect 2200 3220 2220 6380
rect 2480 3220 2500 6380
rect 2200 3200 2500 3220
rect 2910 6380 2990 6500
rect 2910 3220 2920 6380
rect 2980 3220 2990 6380
rect 2910 3210 2990 3220
rect 3010 6380 3090 6390
rect 3010 3220 3020 6380
rect 3080 3220 3090 6380
rect 3010 3210 3090 3220
rect 3110 6380 3190 6500
rect 3110 3220 3120 6380
rect 3180 3220 3190 6380
rect 3110 3210 3190 3220
rect 3610 6380 3690 6390
rect 3610 3220 3620 6380
rect 3680 3220 3690 6380
rect 3610 3100 3690 3220
rect 4110 6380 4190 6390
rect 4110 3220 4120 6380
rect 4180 3220 4190 6380
rect 4110 3100 4190 3220
rect 4610 6380 4690 6390
rect 4610 3220 4620 6380
rect 4680 3220 4690 6380
rect 4610 3100 4690 3220
rect 5110 6380 5190 6500
rect 5110 3220 5120 6380
rect 5180 3220 5190 6380
rect 5110 3210 5190 3220
rect 5210 6380 5290 6390
rect 5210 3220 5220 6380
rect 5280 3220 5290 6380
rect 5210 3210 5290 3220
rect 5310 6380 5390 6500
rect 5310 3220 5320 6380
rect 5380 3220 5390 6380
rect 5310 3210 5390 3220
rect 5810 6380 5890 6500
rect 5810 3220 5820 6380
rect 5880 3220 5890 6380
rect 5810 3210 5890 3220
rect 5910 6380 5990 6390
rect 5910 3220 5920 6380
rect 5980 3220 5990 6380
rect 5910 3210 5990 3220
rect -200 3050 1300 3100
rect -200 2950 -150 3050
rect -50 2950 250 3050
rect 350 2950 750 3050
rect 850 2950 1150 3050
rect 1250 2950 1300 3050
rect -200 2900 1300 2950
rect 3400 3050 4900 3100
rect 3400 2950 3450 3050
rect 3550 2950 3850 3050
rect 3950 2950 4350 3050
rect 4450 2950 4750 3050
rect 4850 2950 4900 3050
rect 3400 2900 4900 2950
<< viali >>
rect -580 7120 -520 10280
rect 2120 7120 2180 10280
rect 4820 7120 4880 10280
rect -1280 3220 -1220 6380
rect -580 3220 -520 6380
rect 1620 3220 1680 6380
rect 2220 3220 2480 6380
rect 3020 3220 3080 6380
rect 5220 3220 5280 6380
rect 5920 3220 5980 6380
<< metal1 >>
rect -1400 10280 6100 10300
rect -1400 7120 -580 10280
rect -520 7120 2120 10280
rect 2180 7120 4820 10280
rect 4880 7120 6100 10280
rect -1400 7100 6100 7120
rect -1400 6380 6100 6400
rect -1400 3220 -1280 6380
rect -1220 3220 -580 6380
rect -520 3220 1620 6380
rect 1680 3220 2220 6380
rect 2480 3220 3020 6380
rect 3080 3220 5220 6380
rect 5280 3220 5920 6380
rect 5980 3220 6100 6380
rect -1400 3200 6100 3220
<< labels >>
flabel metal1 -1400 8600 -1395 8605 0 FreeSans 800 0 0 0 VP
port 1 nsew
flabel metal1 -1400 4600 -1395 4605 0 FreeSans 800 0 0 0 VN
port 2 nsew
flabel poly -1400 10450 -1400 10450 0 FreeSans 800 0 0 0 VBP
port 3 nsew
flabel locali -1400 6750 -1400 6750 0 FreeSans 800 0 0 0 VCN
port 4 nsew
<< end >>
