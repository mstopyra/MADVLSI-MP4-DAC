* NGSPICE file created from first_current_mirror.ext - technology: sky130A

X0 a_2400_28600# a_2400_28600# a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X1 VP VBP a_6000_21500# VP sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X2 a_n200_n400# a_2400_n600# VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=144 ps=41 w=32 l=4
X3 a_n200_29000# a_2400_28600# a_2400_28600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X4 I_OUT I_IN a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X5 a_n200_29000# I_IN I_OUT VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X6 a_n200_29000# VN VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X7 a_2400_n600# VBP a_6000_14300# VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=48 ps=35 w=32 l=4
X8 a_2400_28600# a_2400_28600# a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X9 a_n200_n400# a_2400_n600# a_2400_n600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X10 a_n200_29000# a_2400_28600# a_2400_28600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X11 a_2400_n600# VP VP VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X12 a_2400_n600# a_2400_n600# a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X13 a_n200_29000# a_2400_n600# VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=144 ps=41 w=32 l=4
X14 a_2400_28600# a_2400_28600# a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X15 a_n200_n400# a_2400_n600# a_2400_n600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X16 a_6000_14300# VBP VP VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X17 VP VBP a_6000_14300# VP sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X18 a_n200_n400# a_2400_n600# a_2400_n600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X19 a_2400_n600# a_2400_n600# a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X20 a_2400_28600# a_2400_28600# a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X21 a_n200_n400# I_IN I_IN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X22 I_IN I_IN a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X23 a_6000_21500# VBP a_2400_28600# VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=48 ps=35 w=32 l=4
X24 a_2400_n600# a_2400_n600# a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X25 a_2400_28600# VBP a_6000_21500# VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=48 ps=35 w=32 l=4
X26 a_n200_n400# VN VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X27 VN VN a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X28 VN a_2400_n600# a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=144 pd=41 as=96 ps=70 w=32 l=4
X29 VP VP a_2400_n600# VP sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X30 a_n200_n400# VN VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X31 a_n200_29000# a_2400_28600# a_2400_28600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X32 a_6000_21500# VBP VP VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X33 a_2400_n600# a_2400_n600# a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X34 VN a_2400_n600# a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=144 pd=41 as=96 ps=70 w=32 l=4
X35 a_6000_14300# VBP a_2400_n600# VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=48 ps=35 w=32 l=4
X36 a_n200_29000# VN VN VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X37 VN VN a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X38 VN VN a_n200_n400# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
X39 a_2400_28600# VP VP VP sky130_fd_pr__nfet_01v8 ad=48 pd=35 as=96 ps=70 w=32 l=4
X40 a_n200_n400# a_2400_n600# a_2400_n600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X41 a_n200_29000# a_2400_28600# a_2400_28600# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X42 VP VP a_2400_28600# VP sky130_fd_pr__nfet_01v8 ad=96 pd=70 as=48 ps=35 w=32 l=4
X43 VN VN a_n200_29000# VN sky130_fd_pr__pfet_01v8 ad=96 pd=70 as=96 ps=70 w=32 l=4
.end

